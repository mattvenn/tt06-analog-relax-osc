* NGSPICE file created from osc_parax.ext - technology: sky130A

.subckt osc_parax osc_out VSS VDD
X0 osc_out.t11 osc_a VDD.t27 VDD.t26 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X1 osc_out.t13 osc_a VSS.t17 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X2 osc_out.t10 osc_a VDD.t25 VDD.t24 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X3 VDD osc_a VSS.t18 sky130_fd_pr__res_high_po_0p35 l=18
X4 osc_out.t9 osc_a VDD.t23 VDD.t22 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X5 VDD.t1 osc_b osc_b VDD.t0 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=5.8 ps=40.58 w=20 l=2
**devattr s=232000,8116 d=232000,8116
X6 VDD osc_b VSS.t19 sky130_fd_pr__res_high_po_0p35 l=18
X7 left_cap.t7 right_cap.t5 sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X8 VDD.t21 osc_a osc_out.t8 VDD.t20 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X9 VSS.t26 cset right_cap.t6 VSS.t25 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=20 l=2
**devattr s=232000,8116 d=232000,8116
X10 left_cap.t7 right_cap.t4 sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X11 VDD.t19 osc_a osc_out.t7 VDD.t18 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X12 osc_out.t16 osc_a VSS.t15 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X13 left_cap.t7 right_cap.t3 sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X14 osc_a osc_a VDD.t17 VDD.t16 sky130_fd_pr__pfet_01v8 ad=5.8 pd=40.58 as=0 ps=0 w=20 l=2
**devattr s=232000,8116 d=232000,8116
X15 VDD.t15 osc_a osc_out.t6 VDD.t14 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X16 osc_out.t14 osc_a VSS.t13 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=4452,274 d=2352,140
X17 right_cap.t7 left_cap.t6 sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X18 osc_a osc_b left_cap.t0 VSS.t0 sky130_fd_pr__nfet_01v8 ad=5.8 pd=40.58 as=0 ps=0 w=20 l=2
**devattr s=232000,8116 d=232000,8116
X19 VDD cset VSS.t20 sky130_fd_pr__res_high_po_0p35 l=20
X20 VDD.t5 osc_a osc_out.t5 VDD.t4 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X21 VSS.t11 osc_a osc_out.t17 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X22 right_cap.t8 left_cap.t1 sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X23 right_cap.t7 left_cap.t5 sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X24 left_cap.t7 right_cap.t2 sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X25 VDD.t13 osc_a osc_out.t4 VDD.t12 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X26 left_cap.t2 cset VSS.t24 VSS.t23 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=20 l=2
**devattr s=232000,8116 d=232000,8116
X27 VDD.t7 osc_a osc_out.t3 VDD.t6 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5400,254 d=5500,255
X28 osc_out.t2 osc_a VDD.t11 VDD.t10 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5500,255 d=5400,254
X29 VSS.t9 osc_a osc_out.t12 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X30 VSS.t7 osc_a osc_out.t18 VSS.t6 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=4452,274
X31 right_cap.t7 left_cap.t4 sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X32 VSS.t22 cset cset VSS.t21 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=5.8 ps=40.58 w=20 l=2
**devattr s=232000,8116 d=232000,8116
X33 right_cap.t7 left_cap.t3 sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X34 VSS.t5 osc_a osc_out.t15 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X35 right_cap.t0 osc_a osc_b VSS.t3 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=5.8 ps=40.58 w=20 l=2
**devattr s=232000,8116 d=232000,8116
X36 osc_out.t1 osc_a VDD.t9 VDD.t8 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X37 left_cap.t7 right_cap.t1 sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X38 osc_out.t19 osc_a VSS.t2 VSS.t1 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X39 osc_out.t0 osc_a VDD.t3 VDD.t2 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5400,254 d=5400,254
R0 VDD.n45 VDD.n43 8795.29
R1 VDD.n48 VDD.n47 8795.29
R2 VDD.n37 VDD.n36 8795.29
R3 VDD.n34 VDD.n32 8795.29
R4 VDD.n44 VDD.n40 938.165
R5 VDD.n44 VDD.n41 938.165
R6 VDD.n49 VDD.n41 938.165
R7 VDD.n33 VDD.n29 938.165
R8 VDD.n33 VDD.n30 938.165
R9 VDD.n38 VDD.n30 938.165
R10 VDD.n50 VDD.n49 603.86
R11 VDD.n39 VDD.n38 603.86
R12 VDD.n27 VDD 438.041
R13 VDD.n11 VDD.t13 349.707
R14 VDD.n26 VDD.t27 343.652
R15 VDD.n50 VDD.n40 321.507
R16 VDD.n39 VDD.n29 321.507
R17 VDD.n6 VDD.n5 318.558
R18 VDD.n10 VDD.n9 318.038
R19 VDD.n14 VDD.n8 317.538
R20 VDD.n2 VDD.n1 317.058
R21 VDD.n20 VDD.n4 317.058
R22 VDD.t6 VDD.t10 251.559
R23 VDD.t2 VDD.t12 248.599
R24 VDD.t14 VDD.t2 248.599
R25 VDD.t24 VDD.t14 248.599
R26 VDD.t4 VDD.t24 248.599
R27 VDD.t22 VDD.t4 248.599
R28 VDD.t20 VDD.t22 248.599
R29 VDD.t8 VDD.t20 248.599
R30 VDD.t18 VDD.t8 248.599
R31 VDD.t10 VDD.t18 248.599
R32 VDD.t26 VDD.t6 248.599
R33 VDD VDD.t26 189.409
R34 VDD.n46 VDD.n45 75.6006
R35 VDD.n48 VDD.n42 75.6006
R36 VDD.n37 VDD.n31 75.6006
R37 VDD.n35 VDD.n34 75.6006
R38 VDD.n16 VDD.n15 34.6358
R39 VDD.n20 VDD.n19 34.2593
R40 VDD.n13 VDD.n10 32.7534
R41 VDD.n21 VDD.n2 28.2358
R42 VDD.n1 VDD.t7 27.5805
R43 VDD.n1 VDD.t11 26.5955
R44 VDD.n4 VDD.t9 26.5955
R45 VDD.n4 VDD.t19 26.5955
R46 VDD.n5 VDD.t23 26.5955
R47 VDD.n5 VDD.t21 26.5955
R48 VDD.n8 VDD.t25 26.5955
R49 VDD.n8 VDD.t5 26.5955
R50 VDD.n9 VDD.t3 26.5955
R51 VDD.n9 VDD.t15 26.5955
R52 VDD.n43 VDD.n40 23.1255
R53 VDD.n47 VDD.n41 23.1255
R54 VDD.n32 VDD.n29 23.1255
R55 VDD.n36 VDD.n30 23.1255
R56 VDD.n43 VDD.n42 22.8671
R57 VDD.n47 VDD.n46 22.8671
R58 VDD.n32 VDD.n31 22.8671
R59 VDD.n36 VDD.n35 22.8671
R60 VDD.n26 VDD.n25 22.2123
R61 VDD.n25 VDD.n2 21.4593
R62 VDD.n54 VDD.t1 18.4534
R63 VDD.n51 VDD.t17 18.3784
R64 VDD.n27 VDD.n26 16.5652
R65 VDD.n21 VDD.n20 15.4358
R66 VDD.n14 VDD.n13 12.0476
R67 VDD.n52 VDD.n50 11.113
R68 VDD.n53 VDD.n39 11.113
R69 VDD.n19 VDD.n6 10.1652
R70 VDD.n13 VDD.n12 9.3005
R71 VDD.n15 VDD.n7 9.3005
R72 VDD.n17 VDD.n16 9.3005
R73 VDD.n19 VDD.n18 9.3005
R74 VDD.n20 VDD.n3 9.3005
R75 VDD.n22 VDD.n21 9.3005
R76 VDD.n23 VDD.n2 9.3005
R77 VDD.n25 VDD.n24 9.3005
R78 VDD.n26 VDD.n0 9.3005
R79 VDD.n28 VDD.n27 9.3005
R80 VDD.n11 VDD.n10 6.33664
R81 VDD.n16 VDD.n6 6.02403
R82 VDD.n15 VDD.n14 3.38874
R83 VDD.n45 VDD.n44 3.03329
R84 VDD.n49 VDD.n48 3.03329
R85 VDD.n34 VDD.n33 3.03329
R86 VDD.n38 VDD.n37 3.03329
R87 VDD VDD.n54 1.71914
R88 VDD.n51 VDD 0.586214
R89 VDD.n12 VDD.n11 0.479734
R90 VDD.t16 VDD.n42 0.19977
R91 VDD.n46 VDD.t16 0.19977
R92 VDD.n35 VDD.t0 0.19977
R93 VDD.t0 VDD.n31 0.19977
R94 VDD.n53 VDD.n52 0.118357
R95 VDD.n54 VDD.n53 0.0790714
R96 VDD.n52 VDD.n51 0.0755
R97 VDD.n12 VDD.n7 0.0364375
R98 VDD.n17 VDD.n7 0.0364375
R99 VDD.n18 VDD.n17 0.0364375
R100 VDD.n18 VDD.n3 0.0364375
R101 VDD.n22 VDD.n3 0.0364375
R102 VDD.n23 VDD.n22 0.0364375
R103 VDD.n24 VDD.n23 0.0364375
R104 VDD.n24 VDD.n0 0.0364375
R105 VDD.n28 VDD 0.0184687
R106 VDD VDD.n28 0.009875
R107 VDD.n0 VDD 0.00675
R108 osc_out.n9 osc_out.n8 317.498
R109 osc_out.n11 osc_out.n10 313.452
R110 osc_out.n19 osc_out.n18 313.452
R111 osc_out.n15 osc_out.n14 313.026
R112 osc_out.n13 osc_out.n12 312.618
R113 osc_out.n17 osc_out.n16 312.226
R114 osc_out.n1 osc_out.n0 207.569
R115 osc_out.n3 osc_out.n2 207.569
R116 osc_out.n5 osc_out.n4 207.569
R117 osc_out.n7 osc_out.n6 207.569
R118 osc_out.n9 osc_out.n7 172.8
R119 osc_out.n21 osc_out.n1 60.6123
R120 osc_out.n20 osc_out 57.8991
R121 osc_out.n3 osc_out.n1 50.4476
R122 osc_out.n5 osc_out.n3 50.4476
R123 osc_out.n7 osc_out.n5 50.4476
R124 osc_out.n11 osc_out.n9 45.177
R125 osc_out.n13 osc_out.n11 45.177
R126 osc_out.n17 osc_out.n15 44.8005
R127 osc_out.n19 osc_out.n17 44.424
R128 osc_out.n15 osc_out.n13 44.0476
R129 osc_out.n0 osc_out.t18 40.0005
R130 osc_out.n0 osc_out.t19 40.0005
R131 osc_out.n2 osc_out.t15 40.0005
R132 osc_out.n2 osc_out.t13 40.0005
R133 osc_out.n4 osc_out.t12 40.0005
R134 osc_out.n4 osc_out.t16 40.0005
R135 osc_out.n6 osc_out.t17 40.0005
R136 osc_out.n6 osc_out.t14 40.0005
R137 osc_out.n8 osc_out.t3 26.5955
R138 osc_out.n8 osc_out.t11 26.5955
R139 osc_out.n10 osc_out.t7 26.5955
R140 osc_out.n10 osc_out.t2 26.5955
R141 osc_out.n12 osc_out.t8 26.5955
R142 osc_out.n12 osc_out.t1 26.5955
R143 osc_out.n14 osc_out.t5 26.5955
R144 osc_out.n14 osc_out.t9 26.5955
R145 osc_out.n16 osc_out.t6 26.5955
R146 osc_out.n16 osc_out.t10 26.5955
R147 osc_out.n18 osc_out.t4 26.5955
R148 osc_out.n18 osc_out.t0 26.5955
R149 osc_out.n21 osc_out 12.6066
R150 osc_out osc_out.n19 11.7852
R151 osc_out.n20 osc_out 11.055
R152 osc_out osc_out.n20 2.13383
R153 osc_out osc_out.n21 0.582318
R154 VSS.n83 VSS.n31 16164.9
R155 VSS.n52 VSS.n44 15412.4
R156 VSS.n48 VSS.n44 15412.4
R157 VSS.n52 VSS.n45 15412.4
R158 VSS.n59 VSS.n41 14386.8
R159 VSS.n55 VSS.n41 14386.8
R160 VSS.n59 VSS.n42 14386.8
R161 VSS.n55 VSS.n42 14386.8
R162 VSS.n66 VSS.n38 14386.8
R163 VSS.n62 VSS.n38 14386.8
R164 VSS.n66 VSS.n39 14386.8
R165 VSS.n62 VSS.n39 14386.8
R166 VSS.n74 VSS.n35 14386.8
R167 VSS.n70 VSS.n35 14386.8
R168 VSS.n74 VSS.n36 14386.8
R169 VSS.n70 VSS.n36 14386.8
R170 VSS.n96 VSS.n91 14386.8
R171 VSS.n91 VSS.n27 14386.8
R172 VSS.n27 VSS.n25 14386.8
R173 VSS.n96 VSS.n25 14386.8
R174 VSS.n100 VSS.n21 14386.8
R175 VSS.n100 VSS.n22 14386.8
R176 VSS.n104 VSS.n22 14386.8
R177 VSS.n104 VSS.n21 14386.8
R178 VSS.n81 VSS.n32 14253.5
R179 VSS.n77 VSS.n32 14253.5
R180 VSS.n81 VSS.n33 14253.5
R181 VSS.n77 VSS.n33 14253.5
R182 VSS.n89 VSS.n28 14253.5
R183 VSS.n85 VSS.n28 14253.5
R184 VSS.n89 VSS.n29 14253.5
R185 VSS.n85 VSS.n29 14253.5
R186 VSS.t25 VSS.t6 7681.21
R187 VSS.n84 VSS.n83 4061.27
R188 VSS.n83 VSS.n82 3715.75
R189 VSS.n106 VSS.n105 2820.61
R190 VSS.t19 VSS.n26 2743.15
R191 VSS.n99 VSS.n98 2423.87
R192 VSS.t3 VSS.n90 1780.1
R193 VSS.n98 VSS.t25 1757.41
R194 VSS.n107 VSS.n106 1198.25
R195 VSS.n51 VSS.n46 1001.41
R196 VSS.n49 VSS.n46 1001.41
R197 VSS.n51 VSS.n50 1001.41
R198 VSS.n50 VSS.n49 1001.41
R199 VSS.n58 VSS.n43 934.777
R200 VSS.n56 VSS.n43 934.777
R201 VSS.n58 VSS.n57 934.777
R202 VSS.n57 VSS.n56 934.777
R203 VSS.n65 VSS.n40 934.777
R204 VSS.n63 VSS.n40 934.777
R205 VSS.n65 VSS.n64 934.777
R206 VSS.n64 VSS.n63 934.777
R207 VSS.n73 VSS.n37 934.777
R208 VSS.n71 VSS.n37 934.777
R209 VSS.n73 VSS.n72 934.777
R210 VSS.n72 VSS.n71 934.777
R211 VSS.n95 VSS.n94 934.777
R212 VSS.n94 VSS.n93 934.777
R213 VSS.n93 VSS.n92 934.777
R214 VSS.n95 VSS.n92 934.777
R215 VSS.n101 VSS.n23 934.777
R216 VSS.n102 VSS.n101 934.777
R217 VSS.n103 VSS.n102 934.777
R218 VSS.n103 VSS.n23 934.777
R219 VSS.n80 VSS.n34 926.119
R220 VSS.n78 VSS.n34 926.119
R221 VSS.n80 VSS.n79 926.119
R222 VSS.n79 VSS.n78 926.119
R223 VSS.n88 VSS.n30 926.119
R224 VSS.n86 VSS.n30 926.119
R225 VSS.n88 VSS.n87 926.119
R226 VSS.n87 VSS.n86 926.119
R227 VSS.n76 VSS.n75 903.375
R228 VSS.n61 VSS.n60 903.375
R229 VSS.n31 VSS.n24 807.235
R230 VSS.n68 VSS.n31 685.96
R231 VSS.n105 VSS.t25 648.004
R232 VSS.t3 VSS.n26 648.004
R233 VSS.n69 VSS.n68 586.438
R234 VSS.n99 VSS.n24 553.543
R235 VSS.t12 VSS 477.974
R236 VSS.n54 VSS.n53 346.5
R237 VSS.n68 VSS.n67 316.938
R238 VSS.n30 VSS.n28 292.5
R239 VSS.n28 VSS.t19 292.5
R240 VSS.n79 VSS.n33 292.5
R241 VSS.n33 VSS.t18 292.5
R242 VSS.n34 VSS.n32 292.5
R243 VSS.n32 VSS.t18 292.5
R244 VSS.n50 VSS.n45 292.5
R245 VSS.n46 VSS.n44 292.5
R246 VSS.n44 VSS.t20 292.5
R247 VSS.n87 VSS.n29 292.5
R248 VSS.n29 VSS.t19 292.5
R249 VSS.n47 VSS.n45 285.058
R250 VSS.n5 VSS.t7 245.403
R251 VSS.n16 VSS.t13 240.127
R252 VSS.n97 VSS.t3 235.814
R253 VSS.n75 VSS.t0 235.812
R254 VSS.n69 VSS.t0 235.812
R255 VSS.n67 VSS.t23 235.812
R256 VSS.n61 VSS.t23 235.812
R257 VSS.n60 VSS.t21 235.812
R258 VSS.n54 VSS.t21 235.812
R259 VSS.n7 VSS.n6 200.127
R260 VSS.n10 VSS.n9 200.127
R261 VSS.n14 VSS.n3 200.127
R262 VSS.n97 VSS.n25 175.472
R263 VSS.t6 VSS.t1 162.474
R264 VSS.t1 VSS.t4 162.474
R265 VSS.t4 VSS.t16 162.474
R266 VSS.t16 VSS.t8 162.474
R267 VSS.t8 VSS.t14 162.474
R268 VSS.t14 VSS.t10 162.474
R269 VSS.t10 VSS.t12 162.474
R270 VSS.n90 VSS.t19 159.962
R271 VSS.n84 VSS.t19 159.962
R272 VSS.n98 VSS.n97 158.814
R273 VSS.n106 VSS 143.582
R274 VSS.n48 VSS.n47 107.081
R275 VSS.n82 VSS.t18 101.751
R276 VSS.n76 VSS.t18 101.751
R277 VSS.n53 VSS.t20 101.751
R278 VSS.n24 VSS.t25 94.4616
R279 VSS.n23 VSS.n21 73.1255
R280 VSS.n21 VSS.t25 73.1255
R281 VSS.n96 VSS.n95 73.1255
R282 VSS.t3 VSS.n96 73.1255
R283 VSS.n72 VSS.n36 73.1255
R284 VSS.n36 VSS.t0 73.1255
R285 VSS.n37 VSS.n35 73.1255
R286 VSS.n35 VSS.t0 73.1255
R287 VSS.n64 VSS.n39 73.1255
R288 VSS.n39 VSS.t23 73.1255
R289 VSS.n40 VSS.n38 73.1255
R290 VSS.n38 VSS.t23 73.1255
R291 VSS.n57 VSS.n42 73.1255
R292 VSS.n42 VSS.t21 73.1255
R293 VSS.n43 VSS.n41 73.1255
R294 VSS.n41 VSS.t21 73.1255
R295 VSS.n102 VSS.n22 73.1255
R296 VSS.n22 VSS.t25 73.1255
R297 VSS.n93 VSS.n27 73.1255
R298 VSS.t3 VSS.n27 73.1255
R299 VSS.n6 VSS.t2 40.0005
R300 VSS.n6 VSS.t5 40.0005
R301 VSS.n9 VSS.t17 40.0005
R302 VSS.n9 VSS.t9 40.0005
R303 VSS.n3 VSS.t15 40.0005
R304 VSS.n3 VSS.t11 40.0005
R305 VSS.n20 VSS.n0 34.6358
R306 VSS.n10 VSS.n8 27.4829
R307 VSS.n16 VSS.n0 25.977
R308 VSS.n107 VSS.n20 23.7181
R309 VSS.n14 VSS.n2 22.9652
R310 VSS.n15 VSS.n14 21.4593
R311 VSS.n16 VSS.n15 18.4476
R312 VSS.n10 VSS.n2 16.9417
R313 VSS.n8 VSS.n7 12.424
R314 VSS.n71 VSS.n70 9.59066
R315 VSS.n70 VSS.n69 9.59066
R316 VSS.n74 VSS.n73 9.59066
R317 VSS.n75 VSS.n74 9.59066
R318 VSS.n63 VSS.n62 9.59066
R319 VSS.n62 VSS.n61 9.59066
R320 VSS.n66 VSS.n65 9.59066
R321 VSS.n67 VSS.n66 9.59066
R322 VSS.n56 VSS.n55 9.59066
R323 VSS.n55 VSS.n54 9.59066
R324 VSS.n59 VSS.n58 9.59066
R325 VSS.n60 VSS.n59 9.59066
R326 VSS.n101 VSS.n100 9.59066
R327 VSS.n100 VSS.n99 9.59066
R328 VSS.n104 VSS.n103 9.59066
R329 VSS.n105 VSS.n104 9.59066
R330 VSS.n94 VSS.n91 9.59066
R331 VSS.n91 VSS.n26 9.59066
R332 VSS.n92 VSS.n25 9.59066
R333 VSS.n108 VSS.n107 9.3005
R334 VSS.n8 VSS.n4 9.3005
R335 VSS.n11 VSS.n10 9.3005
R336 VSS.n12 VSS.n2 9.3005
R337 VSS.n14 VSS.n13 9.3005
R338 VSS.n15 VSS.n1 9.3005
R339 VSS.n17 VSS.n16 9.3005
R340 VSS.n18 VSS.n0 9.3005
R341 VSS.n20 VSS.n19 9.3005
R342 VSS.n86 VSS.n85 8.86414
R343 VSS.n85 VSS.n84 8.86414
R344 VSS.n89 VSS.n88 8.86414
R345 VSS.n90 VSS.n89 8.86414
R346 VSS.n78 VSS.n77 8.86414
R347 VSS.n77 VSS.n76 8.86414
R348 VSS.n81 VSS.n80 8.86414
R349 VSS.n82 VSS.n81 8.86414
R350 VSS.n49 VSS.n48 8.1255
R351 VSS.n52 VSS.n51 8.1255
R352 VSS.n53 VSS.n52 8.1255
R353 VSS.n109 VSS.t22 7.61045
R354 VSS.n109 VSS.t24 7.5917
R355 VSS.n111 VSS.t26 7.23714
R356 VSS.n7 VSS.n5 6.81933
R357 VSS.n111 VSS.n110 2.3321
R358 VSS.n47 VSS.t20 2.03318
R359 VSS.n5 VSS.n4 0.688483
R360 VSS.n110 VSS.n109 0.633312
R361 VSS VSS.n111 0.620031
R362 VSS.n110 VSS 0.157907
R363 VSS.n11 VSS.n4 0.0310851
R364 VSS.n12 VSS.n11 0.0310851
R365 VSS.n13 VSS.n12 0.0310851
R366 VSS.n13 VSS.n1 0.0310851
R367 VSS.n17 VSS.n1 0.0310851
R368 VSS.n18 VSS.n17 0.0310851
R369 VSS.n19 VSS.n18 0.0310851
R370 VSS.n108 VSS 0.0157926
R371 VSS VSS.n108 0.00881117
R372 VSS.n19 VSS 0.00581915
R373 left_cap.n1 left_cap.t2 9.38826
R374 left_cap.n1 left_cap.t0 9.20909
R375 left_cap left_cap.n0 7.91907
R376 left_cap left_cap.n1 7.80107
R377 left_cap.n0 left_cap.t1 6.28228
R378 left_cap.t6 left_cap.t4 2.92748
R379 left_cap.t1 left_cap.t3 2.85665
R380 left_cap.t3 left_cap.t5 2.85665
R381 left_cap.t5 left_cap.t6 2.85665
R382 left_cap.n0 left_cap.t7 0.93824
R383 right_cap.n0 right_cap.t6 9.48011
R384 right_cap.n0 right_cap.t0 9.43427
R385 right_cap right_cap.n0 8.02607
R386 right_cap right_cap.t8 7.45138
R387 right_cap.t8 right_cap.t1 3.21837
R388 right_cap.t5 right_cap.t2 2.92748
R389 right_cap.t1 right_cap.t4 2.85665
R390 right_cap.t4 right_cap.t3 2.85665
R391 right_cap.t3 right_cap.t5 2.85665
R392 right_cap.t8 right_cap.t7 1.02493
C0 osc_a left_cap 0.615488f
C1 VDD osc_out 1.21047f
C2 osc_a cset 1.10628f
C3 osc_a right_cap 0.732557f
C4 osc_a VDD 6.18873f
C5 cset left_cap 0.733616f
C6 right_cap left_cap 0.798551p
C7 osc_a osc_b 2.2743f
C8 VDD left_cap 0.063197f
C9 cset right_cap 0.732846f
C10 osc_b left_cap 0.74314f
C11 VDD cset 1.83901f
C12 VDD right_cap 0.07197f
C13 osc_a osc_out 1.4074f
C14 osc_b cset 0.550344f
C15 osc_b right_cap 0.616311f
C16 VDD osc_b 4.08243f
C17 osc_out VSS 2.89777f
C18 VDD VSS 58.746506f
C19 right_cap VSS 93.06754f
C20 osc_a VSS 14.545099f
C21 osc_b VSS 10.9295f
C22 left_cap VSS 0.101902p
C23 cset VSS 17.3869f
C24 right_cap.t7 VSS 0.284166p
C25 right_cap.t8 VSS 0.227929p
C26 right_cap.t2 VSS 56.5149f
C27 right_cap.t5 VSS 56.817f
C28 right_cap.t3 VSS 56.666f
C29 right_cap.t4 VSS 56.666f
C30 right_cap.t1 VSS 56.7594f
C31 right_cap.t6 VSS 0.536933f
C32 right_cap.t0 VSS 0.535327f
C33 right_cap.n0 VSS 1.2457f
C34 left_cap.t7 VSS 0.362111p
C35 left_cap.n0 VSS 0.149859p
C36 left_cap.t4 VSS 56.4468f
C37 left_cap.t6 VSS 56.7485f
C38 left_cap.t5 VSS 56.5977f
C39 left_cap.t3 VSS 56.5977f
C40 left_cap.t1 VSS 57.1758f
C41 left_cap.t0 VSS 0.526352f
C42 left_cap.t2 VSS 0.533095f
C43 left_cap.n1 VSS 1.19422f
C44 VDD.t12 VSS 0.023731f
C45 VDD.t2 VSS 0.007756f
C46 VDD.t14 VSS 0.007756f
C47 VDD.t24 VSS 0.007756f
C48 VDD.t4 VSS 0.007756f
C49 VDD.t22 VSS 0.007756f
C50 VDD.t20 VSS 0.007756f
C51 VDD.t8 VSS 0.007756f
C52 VDD.t18 VSS 0.007756f
C53 VDD.t10 VSS 0.007802f
C54 VDD.t6 VSS 0.007802f
C55 VDD.t26 VSS 0.006833f
C56 VDD.n0 VSS 0.004971f
C57 VDD.t27 VSS 0.002971f
C58 VDD.t11 VSS 7.77e-19
C59 VDD.t7 VSS 8.05e-19
C60 VDD.n1 VSS 0.001746f
C61 VDD.n2 VSS 0.003489f
C62 VDD.n3 VSS 0.008469f
C63 VDD.t9 VSS 7.77e-19
C64 VDD.t19 VSS 7.77e-19
C65 VDD.n4 VSS 0.001717f
C66 VDD.t23 VSS 7.77e-19
C67 VDD.t21 VSS 7.77e-19
C68 VDD.n5 VSS 0.001716f
C69 VDD.n6 VSS 0.00288f
C70 VDD.n7 VSS 0.008469f
C71 VDD.t25 VSS 7.77e-19
C72 VDD.t5 VSS 7.77e-19
C73 VDD.n8 VSS 0.001717f
C74 VDD.t3 VSS 7.77e-19
C75 VDD.t15 VSS 7.77e-19
C76 VDD.n9 VSS 0.001716f
C77 VDD.n10 VSS 0.003521f
C78 VDD.t13 VSS 0.003041f
C79 VDD.n11 VSS 0.01004f
C80 VDD.n12 VSS 0.06337f
C81 VDD.n13 VSS 5.82e-19
C82 VDD.n14 VSS 0.002986f
C83 VDD.n15 VSS 4.94e-19
C84 VDD.n16 VSS 5.28e-19
C85 VDD.n17 VSS 0.008469f
C86 VDD.n18 VSS 0.008469f
C87 VDD.n19 VSS 5.77e-19
C88 VDD.n20 VSS 0.003489f
C89 VDD.n21 VSS 5.67e-19
C90 VDD.n22 VSS 0.008469f
C91 VDD.n23 VSS 0.008469f
C92 VDD.n24 VSS 0.008469f
C93 VDD.n25 VSS 5.67e-19
C94 VDD.n26 VSS 0.003531f
C95 VDD.n27 VSS 0.011317f
C96 VDD.n28 VSS 0.003222f
C97 VDD.t1 VSS 0.083682f
C98 VDD.n29 VSS 0.01661f
C99 VDD.n30 VSS 0.024659f
C100 VDD.n32 VSS 0.024659f
C101 VDD.n33 VSS 0.024418f
C102 VDD.n34 VSS 0.299648f
C103 VDD.t0 VSS 0.460613f
C104 VDD.n36 VSS 0.024659f
C105 VDD.n37 VSS 0.299648f
C106 VDD.n38 VSS 0.020055f
C107 VDD.n39 VSS 0.015426f
C108 VDD.n40 VSS 0.01661f
C109 VDD.n41 VSS 0.024659f
C110 VDD.n43 VSS 0.024659f
C111 VDD.n44 VSS 0.024418f
C112 VDD.n45 VSS 0.299648f
C113 VDD.t16 VSS 0.460613f
C114 VDD.n47 VSS 0.024659f
C115 VDD.n48 VSS 0.299648f
C116 VDD.n49 VSS 0.020055f
C117 VDD.n50 VSS 0.015426f
C118 VDD.t17 VSS 0.093994f
C119 VDD.n51 VSS 1.59338f
C120 VDD.n52 VSS 0.460335f
C121 VDD.n53 VSS 0.46839f
C122 VDD.n54 VSS 2.59477f
.ends

