VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_mattvenn_relax_osc
  CLASS BLOCK ;
  FOREIGN tt_um_mattvenn_relax_osc ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 156.560 0.000 157.160 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 134.480 0.000 135.080 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 112.400 0.000 113.000 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.320 0.000 90.920 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.240 0.000 68.840 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.160 0.000 46.760 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 24.080 0.000 24.680 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 2.000 0.000 2.600 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 49.000 5.000 50.500 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 54.950 186.670 56.960 212.490 ;
        RECT 58.950 186.670 62.910 208.770 ;
        RECT 68.950 186.670 72.910 208.770 ;
        RECT 78.950 186.670 82.910 208.770 ;
        RECT 88.950 186.670 90.960 210.490 ;
      LAYER nwell ;
        RECT 94.950 186.670 98.910 208.860 ;
        RECT 104.950 186.670 108.910 208.860 ;
      LAYER pwell ;
        RECT 112.950 186.670 114.960 210.490 ;
        RECT 120.950 186.670 124.910 208.770 ;
        RECT 131.950 186.670 135.910 208.770 ;
      LAYER nwell ;
        RECT 143.150 198.315 149.510 199.920 ;
      LAYER pwell ;
        RECT 144.285 197.115 148.235 197.795 ;
        RECT 143.490 196.925 143.660 197.095 ;
      LAYER li1 ;
        RECT 55.130 212.140 56.780 212.310 ;
        RECT 55.130 187.020 55.300 212.140 ;
        RECT 55.780 209.500 56.130 211.660 ;
        RECT 55.780 187.500 56.130 189.660 ;
        RECT 56.610 187.020 56.780 212.140 ;
        RECT 89.130 210.140 90.780 210.310 ;
        RECT 55.130 186.850 56.780 187.020 ;
        RECT 59.130 208.420 62.730 208.590 ;
        RECT 59.130 187.020 59.300 208.420 ;
        RECT 59.930 207.910 61.930 208.080 ;
        RECT 59.700 187.700 59.870 207.740 ;
        RECT 61.990 187.700 62.160 207.740 ;
        RECT 59.930 187.360 61.930 187.530 ;
        RECT 62.560 187.020 62.730 208.420 ;
        RECT 59.130 186.850 62.730 187.020 ;
        RECT 69.130 208.420 72.730 208.590 ;
        RECT 69.130 187.020 69.300 208.420 ;
        RECT 69.930 207.910 71.930 208.080 ;
        RECT 69.700 187.700 69.870 207.740 ;
        RECT 71.990 187.700 72.160 207.740 ;
        RECT 69.930 187.360 71.930 187.530 ;
        RECT 72.560 187.020 72.730 208.420 ;
        RECT 69.130 186.850 72.730 187.020 ;
        RECT 79.130 208.420 82.730 208.590 ;
        RECT 79.130 187.020 79.300 208.420 ;
        RECT 79.930 207.910 81.930 208.080 ;
        RECT 79.700 187.700 79.870 207.740 ;
        RECT 81.990 187.700 82.160 207.740 ;
        RECT 79.930 187.360 81.930 187.530 ;
        RECT 82.560 187.020 82.730 208.420 ;
        RECT 79.130 186.850 82.730 187.020 ;
        RECT 89.130 187.020 89.300 210.140 ;
        RECT 89.780 207.500 90.130 209.660 ;
        RECT 89.780 187.500 90.130 189.660 ;
        RECT 90.610 187.020 90.780 210.140 ;
        RECT 113.130 210.140 114.780 210.310 ;
        RECT 89.130 186.850 90.780 187.020 ;
        RECT 95.130 208.510 98.730 208.680 ;
        RECT 95.130 187.020 95.300 208.510 ;
        RECT 95.930 208.000 97.930 208.170 ;
        RECT 95.700 187.745 95.870 207.785 ;
        RECT 97.990 187.745 98.160 207.785 ;
        RECT 98.560 206.040 98.730 208.510 ;
        RECT 105.130 208.510 108.730 208.680 ;
        RECT 105.130 206.040 105.300 208.510 ;
        RECT 105.930 208.000 107.930 208.170 ;
        RECT 98.480 205.700 98.820 206.040 ;
        RECT 105.080 205.700 105.420 206.040 ;
        RECT 95.930 187.360 97.930 187.530 ;
        RECT 98.560 187.020 98.730 205.700 ;
        RECT 95.130 186.850 98.730 187.020 ;
        RECT 105.130 187.020 105.300 205.700 ;
        RECT 105.700 187.745 105.870 207.785 ;
        RECT 107.990 187.745 108.160 207.785 ;
        RECT 105.930 187.360 107.930 187.530 ;
        RECT 108.560 187.020 108.730 208.510 ;
        RECT 105.130 186.850 108.730 187.020 ;
        RECT 113.130 187.020 113.300 210.140 ;
        RECT 113.780 207.500 114.130 209.660 ;
        RECT 113.780 187.500 114.130 189.660 ;
        RECT 114.610 187.020 114.780 210.140 ;
        RECT 113.130 186.850 114.780 187.020 ;
        RECT 121.130 208.420 124.730 208.590 ;
        RECT 121.130 187.020 121.300 208.420 ;
        RECT 121.930 207.910 123.930 208.080 ;
        RECT 121.700 187.700 121.870 207.740 ;
        RECT 123.990 187.700 124.160 207.740 ;
        RECT 121.930 187.360 123.930 187.530 ;
        RECT 124.560 187.020 124.730 208.420 ;
        RECT 121.130 186.850 124.730 187.020 ;
        RECT 132.130 208.420 135.730 208.590 ;
        RECT 132.130 187.020 132.300 208.420 ;
        RECT 132.930 207.910 134.930 208.080 ;
        RECT 132.700 187.700 132.870 207.740 ;
        RECT 134.990 187.700 135.160 207.740 ;
        RECT 132.930 187.360 134.930 187.530 ;
        RECT 135.560 187.020 135.730 208.420 ;
        RECT 143.340 199.645 149.320 199.815 ;
        RECT 143.475 198.810 143.735 199.645 ;
        RECT 143.905 198.640 144.145 199.445 ;
        RECT 144.315 198.810 144.575 199.645 ;
        RECT 144.745 198.640 144.985 199.445 ;
        RECT 145.155 198.810 145.415 199.645 ;
        RECT 145.585 198.640 145.835 199.445 ;
        RECT 146.005 198.810 146.250 199.645 ;
        RECT 146.420 198.640 146.665 199.445 ;
        RECT 146.835 198.810 147.090 199.645 ;
        RECT 147.260 198.640 147.515 199.445 ;
        RECT 147.685 198.810 147.935 199.645 ;
        RECT 148.105 198.640 148.345 199.445 ;
        RECT 148.515 198.810 148.770 199.645 ;
        RECT 143.455 198.570 148.780 198.640 ;
        RECT 143.455 198.470 152.650 198.570 ;
        RECT 143.455 197.875 143.625 198.470 ;
        RECT 143.795 198.045 148.205 198.300 ;
        RECT 148.450 197.875 152.650 198.470 ;
        RECT 143.455 197.770 152.650 197.875 ;
        RECT 143.455 197.705 148.780 197.770 ;
        RECT 144.375 197.095 144.705 197.535 ;
        RECT 144.875 197.290 145.065 197.705 ;
        RECT 145.235 197.095 145.565 197.535 ;
        RECT 145.735 197.290 145.925 197.705 ;
        RECT 146.095 197.095 146.425 197.535 ;
        RECT 146.595 197.290 146.785 197.705 ;
        RECT 146.955 197.095 147.285 197.535 ;
        RECT 147.455 197.290 147.645 197.705 ;
        RECT 147.815 197.095 148.145 197.535 ;
        RECT 143.340 196.925 149.320 197.095 ;
        RECT 132.130 186.850 135.730 187.020 ;
      LAYER mcon ;
        RECT 55.860 209.585 56.050 211.570 ;
        RECT 55.860 187.590 56.050 189.575 ;
        RECT 60.010 207.910 61.850 208.080 ;
        RECT 59.700 187.780 59.870 207.660 ;
        RECT 61.990 187.780 62.160 207.660 ;
        RECT 60.010 187.360 61.850 187.530 ;
        RECT 70.010 207.910 71.850 208.080 ;
        RECT 69.700 187.780 69.870 207.660 ;
        RECT 71.990 187.780 72.160 207.660 ;
        RECT 70.010 187.360 71.850 187.530 ;
        RECT 80.010 207.910 81.850 208.080 ;
        RECT 79.700 187.780 79.870 207.660 ;
        RECT 81.990 187.780 82.160 207.660 ;
        RECT 80.010 187.360 81.850 187.530 ;
        RECT 89.860 207.585 90.050 209.570 ;
        RECT 89.860 187.590 90.050 189.575 ;
        RECT 96.010 208.000 97.850 208.170 ;
        RECT 95.700 187.825 95.870 207.705 ;
        RECT 97.990 187.825 98.160 207.705 ;
        RECT 106.010 208.000 107.850 208.170 ;
        RECT 98.480 205.700 98.820 206.040 ;
        RECT 105.080 205.700 105.420 206.040 ;
        RECT 96.010 187.360 97.850 187.530 ;
        RECT 105.700 187.825 105.870 207.705 ;
        RECT 107.990 187.825 108.160 207.705 ;
        RECT 106.010 187.360 107.850 187.530 ;
        RECT 113.860 207.585 114.050 209.570 ;
        RECT 113.860 187.590 114.050 189.575 ;
        RECT 122.010 207.910 123.850 208.080 ;
        RECT 121.700 187.780 121.870 207.660 ;
        RECT 123.990 187.780 124.160 207.660 ;
        RECT 122.010 187.360 123.850 187.530 ;
        RECT 133.010 207.910 134.850 208.080 ;
        RECT 132.700 187.780 132.870 207.660 ;
        RECT 134.990 187.780 135.160 207.660 ;
        RECT 133.010 187.360 134.850 187.530 ;
        RECT 143.485 199.645 143.655 199.815 ;
        RECT 143.945 199.645 144.115 199.815 ;
        RECT 144.405 199.645 144.575 199.815 ;
        RECT 144.865 199.645 145.035 199.815 ;
        RECT 145.325 199.645 145.495 199.815 ;
        RECT 145.785 199.645 145.955 199.815 ;
        RECT 146.245 199.645 146.415 199.815 ;
        RECT 146.705 199.645 146.875 199.815 ;
        RECT 147.165 199.645 147.335 199.815 ;
        RECT 147.625 199.645 147.795 199.815 ;
        RECT 148.085 199.645 148.255 199.815 ;
        RECT 148.545 199.645 148.715 199.815 ;
        RECT 149.005 199.645 149.175 199.815 ;
        RECT 146.765 198.085 146.935 198.255 ;
        RECT 151.880 197.800 152.620 198.540 ;
        RECT 143.485 196.925 143.655 197.095 ;
        RECT 143.945 196.925 144.115 197.095 ;
        RECT 144.405 196.925 144.575 197.095 ;
        RECT 144.865 196.925 145.035 197.095 ;
        RECT 145.325 196.925 145.495 197.095 ;
        RECT 145.785 196.925 145.955 197.095 ;
        RECT 146.245 196.925 146.415 197.095 ;
        RECT 146.705 196.925 146.875 197.095 ;
        RECT 147.165 196.925 147.335 197.095 ;
        RECT 147.625 196.925 147.795 197.095 ;
        RECT 148.085 196.925 148.255 197.095 ;
        RECT 148.545 196.925 148.715 197.095 ;
        RECT 149.005 196.925 149.175 197.095 ;
      LAYER met1 ;
        RECT 58.850 214.270 142.850 218.670 ;
        RECT 55.450 213.470 142.850 214.270 ;
        RECT 55.455 210.875 56.245 213.470 ;
        RECT 58.850 211.670 142.850 213.470 ;
        RECT 89.750 211.175 90.150 211.670 ;
        RECT 55.830 209.525 56.080 210.875 ;
        RECT 57.150 209.270 71.350 210.070 ;
        RECT 57.150 191.670 57.950 209.270 ;
        RECT 70.650 208.110 71.150 209.270 ;
        RECT 80.800 208.110 81.300 209.950 ;
        RECT 59.950 207.880 61.910 208.110 ;
        RECT 69.950 207.880 71.910 208.110 ;
        RECT 79.950 207.880 81.910 208.110 ;
        RECT 89.750 207.970 90.155 211.175 ;
        RECT 59.670 191.670 59.900 207.720 ;
        RECT 61.960 192.070 62.190 207.720 ;
        RECT 69.670 192.070 69.900 207.720 ;
        RECT 70.650 207.570 71.150 207.880 ;
        RECT 71.960 206.170 72.190 207.720 ;
        RECT 76.060 206.170 76.660 206.200 ;
        RECT 79.670 206.170 79.900 207.720 ;
        RECT 80.800 207.420 81.300 207.880 ;
        RECT 71.850 205.570 80.050 206.170 ;
        RECT 57.150 190.870 60.250 191.670 ;
        RECT 55.830 188.670 56.080 189.635 ;
        RECT 57.150 188.670 57.950 190.870 ;
        RECT 55.650 187.870 57.950 188.670 ;
        RECT 55.830 187.530 56.080 187.870 ;
        RECT 57.150 185.570 57.950 187.870 ;
        RECT 59.670 187.720 59.900 190.870 ;
        RECT 61.250 190.470 70.450 192.070 ;
        RECT 60.450 187.560 61.250 187.870 ;
        RECT 61.960 187.720 62.190 190.470 ;
        RECT 59.950 187.330 61.910 187.560 ;
        RECT 60.450 185.570 61.250 187.330 ;
        RECT 57.150 184.770 61.250 185.570 ;
        RECT 65.250 182.370 66.850 190.470 ;
        RECT 69.670 187.720 69.900 190.470 ;
        RECT 71.960 187.720 72.190 205.570 ;
        RECT 76.060 205.540 76.660 205.570 ;
        RECT 79.670 187.720 79.900 205.570 ;
        RECT 81.960 188.820 82.190 207.720 ;
        RECT 89.830 207.525 90.080 207.970 ;
        RECT 94.250 207.070 94.650 211.670 ;
        RECT 95.950 207.970 97.910 208.200 ;
        RECT 95.670 207.070 95.900 207.765 ;
        RECT 94.250 206.670 96.050 207.070 ;
        RECT 89.830 188.820 90.080 189.635 ;
        RECT 81.700 188.320 90.200 188.820 ;
        RECT 81.960 187.720 82.190 188.320 ;
        RECT 69.950 187.330 71.910 187.560 ;
        RECT 79.950 187.330 81.910 187.560 ;
        RECT 87.600 185.970 88.100 188.320 ;
        RECT 89.830 187.530 90.080 188.320 ;
        RECT 95.670 187.765 95.900 206.670 ;
        RECT 97.960 189.120 98.190 207.765 ;
        RECT 98.450 205.640 98.850 211.670 ;
        RECT 105.050 205.640 105.450 211.670 ;
        RECT 105.950 207.970 107.910 208.200 ;
        RECT 103.770 197.720 104.330 198.220 ;
        RECT 99.900 189.120 100.400 195.550 ;
        RECT 97.700 188.620 100.400 189.120 ;
        RECT 97.960 187.765 98.190 188.620 ;
        RECT 96.700 187.560 97.200 187.720 ;
        RECT 95.950 187.330 97.910 187.560 ;
        RECT 96.700 185.970 97.200 187.330 ;
        RECT 99.900 185.970 100.400 188.620 ;
        RECT 103.800 192.740 104.300 197.720 ;
        RECT 103.800 191.940 104.350 192.740 ;
        RECT 103.800 189.120 104.300 191.940 ;
        RECT 105.670 189.120 105.900 207.765 ;
        RECT 107.960 207.070 108.190 207.765 ;
        RECT 109.450 207.070 109.850 211.670 ;
        RECT 113.750 207.470 114.150 211.670 ;
        RECT 119.150 211.640 119.650 211.670 ;
        RECT 122.670 209.420 123.230 209.920 ;
        RECT 122.700 208.110 123.200 209.420 ;
        RECT 133.700 208.110 134.200 209.800 ;
        RECT 121.950 207.880 123.910 208.110 ;
        RECT 132.950 207.880 134.910 208.110 ;
        RECT 107.850 206.670 109.850 207.070 ;
        RECT 107.960 195.740 108.190 206.670 ;
        RECT 107.550 194.940 108.750 195.740 ;
        RECT 103.800 188.620 106.100 189.120 ;
        RECT 103.800 185.970 104.300 188.620 ;
        RECT 105.670 187.765 105.900 188.620 ;
        RECT 107.960 187.765 108.190 194.940 ;
        RECT 113.830 188.920 114.080 189.635 ;
        RECT 113.700 188.820 115.800 188.920 ;
        RECT 121.670 188.820 121.900 207.720 ;
        RECT 122.700 207.520 123.200 207.880 ;
        RECT 133.700 207.720 134.200 207.880 ;
        RECT 123.960 206.270 124.190 207.720 ;
        RECT 128.020 206.270 128.620 206.300 ;
        RECT 132.670 206.270 132.900 207.720 ;
        RECT 123.750 205.670 133.050 206.270 ;
        RECT 113.700 188.420 122.100 188.820 ;
        RECT 105.950 187.330 107.910 187.560 ;
        RECT 113.830 187.530 114.080 188.420 ;
        RECT 115.300 188.320 122.100 188.420 ;
        RECT 106.800 185.970 107.300 187.330 ;
        RECT 115.300 185.970 115.800 188.320 ;
        RECT 121.670 187.720 121.900 188.320 ;
        RECT 123.960 187.720 124.190 205.670 ;
        RECT 128.020 205.640 128.620 205.670 ;
        RECT 132.670 187.720 132.900 205.670 ;
        RECT 134.960 192.570 135.190 207.720 ;
        RECT 137.150 201.070 138.750 211.670 ;
        RECT 137.050 199.470 150.750 201.070 ;
        RECT 140.550 198.270 141.250 198.670 ;
        RECT 152.550 198.570 158.450 200.670 ;
        RECT 146.705 198.270 146.995 198.285 ;
        RECT 140.550 198.070 146.995 198.270 ;
        RECT 140.550 197.770 141.250 198.070 ;
        RECT 146.705 198.055 146.995 198.070 ;
        RECT 151.820 197.770 158.450 198.570 ;
        RECT 143.340 196.970 149.320 197.250 ;
        RECT 136.950 195.370 150.650 196.970 ;
        RECT 136.950 192.570 138.550 195.370 ;
        RECT 152.550 195.070 158.450 197.770 ;
        RECT 134.250 190.970 138.550 192.570 ;
        RECT 134.960 187.720 135.190 190.970 ;
        RECT 121.950 187.330 123.910 187.560 ;
        RECT 132.950 187.330 134.910 187.560 ;
        RECT 87.600 185.470 100.450 185.970 ;
        RECT 103.750 185.470 115.800 185.970 ;
        RECT 136.950 182.370 138.550 190.970 ;
        RECT 57.350 176.970 140.750 182.370 ;
      LAYER via ;
        RECT 70.650 209.270 71.150 209.770 ;
        RECT 80.800 209.420 81.300 209.920 ;
        RECT 76.060 205.570 76.660 206.170 ;
        RECT 103.800 197.720 104.300 198.220 ;
        RECT 99.900 195.020 100.400 195.520 ;
        RECT 122.700 209.420 123.200 209.920 ;
        RECT 133.700 209.270 134.200 209.770 ;
        RECT 128.020 205.670 128.620 206.270 ;
        RECT 140.600 197.920 141.100 198.420 ;
      LAYER met2 ;
        RECT 118.300 210.420 141.200 210.920 ;
        RECT 118.300 209.920 118.800 210.420 ;
        RECT 122.700 209.920 123.200 209.950 ;
        RECT 70.650 209.770 71.150 209.800 ;
        RECT 70.650 209.270 76.345 209.770 ;
        RECT 80.770 209.420 85.800 209.920 ;
        RECT 70.650 209.240 71.150 209.270 ;
        RECT 76.030 205.570 76.690 206.170 ;
        RECT 76.060 173.800 76.660 205.570 ;
        RECT 85.300 198.220 85.800 209.420 ;
        RECT 118.300 209.420 123.200 209.920 ;
        RECT 127.425 209.770 127.875 209.790 ;
        RECT 103.800 198.220 104.300 198.250 ;
        RECT 85.300 197.720 104.300 198.220 ;
        RECT 103.800 197.690 104.300 197.720 ;
        RECT 118.300 195.520 118.800 209.420 ;
        RECT 122.700 209.390 123.200 209.420 ;
        RECT 127.400 209.270 134.340 209.770 ;
        RECT 127.425 209.250 127.875 209.270 ;
        RECT 140.700 208.760 141.200 210.420 ;
        RECT 140.600 207.420 141.200 208.760 ;
        RECT 127.990 205.670 128.650 206.270 ;
        RECT 99.870 195.020 118.800 195.520 ;
        RECT 76.060 173.200 80.255 173.800 ;
        RECT 128.020 172.820 128.620 205.670 ;
        RECT 140.600 197.890 141.100 207.420 ;
        RECT 127.975 172.220 128.665 172.820 ;
      LAYER via2 ;
        RECT 75.800 209.270 76.300 209.770 ;
        RECT 127.425 209.295 127.875 209.745 ;
        RECT 79.610 173.200 80.210 173.800 ;
        RECT 128.020 172.220 128.620 172.820 ;
      LAYER met3 ;
        RECT 75.775 209.770 76.325 209.795 ;
        RECT 75.775 209.270 127.900 209.770 ;
        RECT 75.775 209.245 76.325 209.270 ;
        RECT 79.585 173.800 80.235 173.825 ;
        RECT 79.585 173.200 81.810 173.800 ;
        RECT 79.585 173.175 80.235 173.200 ;
        RECT 127.995 172.820 128.645 172.845 ;
        RECT 123.960 172.220 128.645 172.820 ;
        RECT 127.995 172.195 128.645 172.220 ;
        RECT 69.350 140.610 101.210 171.010 ;
        RECT 105.730 141.190 137.590 171.590 ;
        RECT 69.350 109.010 101.210 139.410 ;
        RECT 105.730 109.590 137.590 139.990 ;
        RECT 69.350 77.410 101.210 107.810 ;
        RECT 105.730 77.990 137.590 108.390 ;
        RECT 69.350 45.810 101.210 76.210 ;
        RECT 105.730 46.390 137.590 76.790 ;
        RECT 69.350 14.210 101.210 44.610 ;
        RECT 105.730 14.790 137.590 45.190 ;
      LAYER via3 ;
        RECT 81.180 173.200 81.780 173.800 ;
        RECT 123.990 172.220 124.590 172.820 ;
        RECT 100.790 140.750 101.110 170.870 ;
        RECT 137.170 141.330 137.490 171.450 ;
        RECT 100.790 109.150 101.110 139.270 ;
        RECT 137.170 109.730 137.490 139.850 ;
        RECT 100.790 77.550 101.110 107.670 ;
        RECT 137.170 78.130 137.490 108.250 ;
        RECT 100.790 45.950 101.110 76.070 ;
        RECT 137.170 46.530 137.490 76.650 ;
        RECT 100.790 14.350 101.110 44.470 ;
        RECT 137.170 14.930 137.490 45.050 ;
      LAYER met4 ;
        RECT 3.990 223.550 4.290 224.760 ;
        RECT 7.670 223.550 7.970 224.760 ;
        RECT 11.350 223.550 11.650 224.760 ;
        RECT 15.030 223.550 15.330 224.760 ;
        RECT 18.710 223.550 19.010 224.760 ;
        RECT 22.390 223.550 22.690 224.760 ;
        RECT 26.070 223.550 26.370 224.760 ;
        RECT 29.750 223.550 30.050 224.760 ;
        RECT 33.430 223.550 33.730 224.760 ;
        RECT 37.110 223.550 37.410 224.760 ;
        RECT 40.790 223.550 41.090 224.760 ;
        RECT 44.470 223.550 44.770 224.760 ;
        RECT 48.150 223.550 48.450 224.760 ;
        RECT 51.830 223.550 52.130 224.760 ;
        RECT 55.510 223.550 55.810 224.760 ;
        RECT 59.190 223.550 59.490 224.760 ;
        RECT 62.870 223.550 63.170 224.760 ;
        RECT 66.550 223.550 66.850 224.760 ;
        RECT 70.230 223.550 70.530 224.760 ;
        RECT 73.910 223.550 74.210 224.760 ;
        RECT 77.590 223.550 77.890 224.760 ;
        RECT 81.270 223.550 81.570 224.760 ;
        RECT 84.950 223.550 85.250 224.760 ;
        RECT 88.630 223.550 88.930 224.760 ;
        RECT 2.760 222.050 89.560 223.550 ;
        RECT 49.000 220.760 50.500 222.050 ;
        RECT 81.175 173.800 81.785 173.805 ;
        RECT 84.290 173.800 137.600 173.870 ;
        RECT 81.175 173.350 137.600 173.800 ;
        RECT 81.175 173.200 85.120 173.350 ;
        RECT 81.175 173.195 81.785 173.200 ;
        RECT 84.290 170.615 84.810 173.200 ;
        RECT 123.985 172.820 124.595 172.825 ;
        RECT 119.240 172.800 124.595 172.820 ;
        RECT 100.610 172.280 124.595 172.800 ;
        RECT 100.610 171.610 101.130 172.280 ;
        RECT 119.240 172.220 124.595 172.280 ;
        RECT 69.745 141.005 99.355 170.615 ;
        RECT 100.610 166.340 101.210 171.610 ;
        RECT 120.670 171.195 121.190 172.220 ;
        RECT 123.985 172.215 124.595 172.220 ;
        RECT 137.080 172.190 137.600 173.350 ;
        RECT 84.290 139.015 84.810 141.005 ;
        RECT 69.745 109.405 99.355 139.015 ;
        RECT 84.290 107.415 84.810 109.405 ;
        RECT 69.745 77.805 99.355 107.415 ;
        RECT 84.290 75.815 84.810 77.805 ;
        RECT 69.745 46.205 99.355 75.815 ;
        RECT 84.290 44.215 84.810 46.205 ;
        RECT 69.745 14.605 99.355 44.215 ;
        RECT 84.290 13.610 84.810 14.605 ;
        RECT 100.690 13.610 101.210 166.340 ;
        RECT 106.125 141.585 135.735 171.195 ;
        RECT 137.070 165.730 137.600 172.190 ;
        RECT 120.670 139.595 121.190 141.585 ;
        RECT 106.125 109.985 135.735 139.595 ;
        RECT 120.670 107.995 121.190 109.985 ;
        RECT 106.125 78.385 135.735 107.995 ;
        RECT 120.670 76.395 121.190 78.385 ;
        RECT 106.125 46.785 135.735 76.395 ;
        RECT 120.670 44.795 121.190 46.785 ;
        RECT 106.125 15.185 135.735 44.795 ;
        RECT 120.670 14.190 121.190 15.185 ;
        RECT 137.070 14.190 137.590 165.730 ;
  END
END tt_um_mattvenn_relax_osc
END LIBRARY

