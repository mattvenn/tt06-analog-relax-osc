** sch_path: /home/matt/work/asic-workshop/shuttle-2404/tt06-analog-relax-osc/xschem/osc.sch
.subckt osc osc_out VDD VSS osc_a
*.PININFO osc_out:B VDD:B VSS:B osc_a:B
XM1 osc_a osc_b left_cap VSS sky130_fd_pr__nfet_01v8 L=2 W=20 nf=1 m=1
XM2 osc_b osc_a right_cap VSS sky130_fd_pr__nfet_01v8 L=2 W=20 nf=1 m=1
XM3 osc_b osc_b VDD VDD sky130_fd_pr__pfet_01v8 L=2 W=20 nf=1 m=1
XM4 osc_a osc_a VDD VDD sky130_fd_pr__pfet_01v8 L=2 W=20 nf=1 m=1
XR1 osc_a VDD VSS sky130_fd_pr__res_high_po_0p35 L=18 mult=1 m=1
XR2 osc_b VDD VSS sky130_fd_pr__res_high_po_0p35 L=18 mult=1 m=1
XC1 right_cap left_cap sky130_fd_pr__cap_mim_m3_1 W=30 L=30 m=5
XM5 cset cset VSS VSS sky130_fd_pr__nfet_01v8 L=2 W=20 nf=1 m=1
XM6 left_cap cset VSS VSS sky130_fd_pr__nfet_01v8 L=2 W=20 nf=1 m=1
XR3 cset VDD VSS sky130_fd_pr__res_high_po_0p35 L=20 mult=1 m=1
XM8 right_cap cset VSS VSS sky130_fd_pr__nfet_01v8 L=2 W=20 nf=1 m=1
x1 osc_a VSS VSS VDD VDD osc_out sky130_fd_sc_hd__clkinv_8
XC2 left_cap right_cap sky130_fd_pr__cap_mim_m3_1 W=30 L=30 m=5
.ends
.end
