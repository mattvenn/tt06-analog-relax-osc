magic
tech sky130A
magscale 1 2
timestamp 1710760421
<< metal3 >>
rect -3186 15652 3186 15680
rect -3186 9628 3102 15652
rect 3166 9628 3186 15652
rect -3186 9600 3186 9628
rect -3186 9332 3186 9360
rect -3186 3308 3102 9332
rect 3166 3308 3186 9332
rect -3186 3280 3186 3308
rect -3186 3012 3186 3040
rect -3186 -3012 3102 3012
rect 3166 -3012 3186 3012
rect -3186 -3040 3186 -3012
rect -3186 -3308 3186 -3280
rect -3186 -9332 3102 -3308
rect 3166 -9332 3186 -3308
rect -3186 -9360 3186 -9332
rect -3186 -9628 3186 -9600
rect -3186 -15652 3102 -9628
rect 3166 -15652 3186 -9628
rect -3186 -15680 3186 -15652
<< via3 >>
rect 3102 9628 3166 15652
rect 3102 3308 3166 9332
rect 3102 -3012 3166 3012
rect 3102 -9332 3166 -3308
rect 3102 -15652 3166 -9628
<< mimcap >>
rect -3146 15600 2854 15640
rect -3146 9680 -3106 15600
rect 2814 9680 2854 15600
rect -3146 9640 2854 9680
rect -3146 9280 2854 9320
rect -3146 3360 -3106 9280
rect 2814 3360 2854 9280
rect -3146 3320 2854 3360
rect -3146 2960 2854 3000
rect -3146 -2960 -3106 2960
rect 2814 -2960 2854 2960
rect -3146 -3000 2854 -2960
rect -3146 -3360 2854 -3320
rect -3146 -9280 -3106 -3360
rect 2814 -9280 2854 -3360
rect -3146 -9320 2854 -9280
rect -3146 -9680 2854 -9640
rect -3146 -15600 -3106 -9680
rect 2814 -15600 2854 -9680
rect -3146 -15640 2854 -15600
<< mimcapcontact >>
rect -3106 9680 2814 15600
rect -3106 3360 2814 9280
rect -3106 -2960 2814 2960
rect -3106 -9280 2814 -3360
rect -3106 -15600 2814 -9680
<< metal4 >>
rect -198 15601 -94 15800
rect 3082 15652 3186 15800
rect -3107 15600 2815 15601
rect -3107 9680 -3106 15600
rect 2814 9680 2815 15600
rect -3107 9679 2815 9680
rect -198 9281 -94 9679
rect 3082 9628 3102 15652
rect 3166 9628 3186 15652
rect 3082 9332 3186 9628
rect -3107 9280 2815 9281
rect -3107 3360 -3106 9280
rect 2814 3360 2815 9280
rect -3107 3359 2815 3360
rect -198 2961 -94 3359
rect 3082 3308 3102 9332
rect 3166 3308 3186 9332
rect 3082 3012 3186 3308
rect -3107 2960 2815 2961
rect -3107 -2960 -3106 2960
rect 2814 -2960 2815 2960
rect -3107 -2961 2815 -2960
rect -198 -3359 -94 -2961
rect 3082 -3012 3102 3012
rect 3166 -3012 3186 3012
rect 3082 -3308 3186 -3012
rect -3107 -3360 2815 -3359
rect -3107 -9280 -3106 -3360
rect 2814 -9280 2815 -3360
rect -3107 -9281 2815 -9280
rect -198 -9679 -94 -9281
rect 3082 -9332 3102 -3308
rect 3166 -9332 3186 -3308
rect 3082 -9628 3186 -9332
rect -3107 -9680 2815 -9679
rect -3107 -15600 -3106 -9680
rect 2814 -15600 2815 -9680
rect -3107 -15601 2815 -15600
rect -198 -15800 -94 -15601
rect 3082 -15652 3102 -9628
rect 3166 -15652 3186 -9628
rect 3082 -15800 3186 -15652
<< properties >>
string FIXED_BBOX -3186 9600 2894 15680
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 30.0 l 30.0 val 1.822k carea 2.00 cperi 0.19 nx 1 ny 5 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
