VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_mattvenn_relax_osc
  CLASS BLOCK ;
  FOREIGN tt_um_mattvenn_relax_osc ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 156.560 0.000 157.160 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 134.480 0.000 135.080 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 112.400 0.000 113.000 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.320 0.000 90.920 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.240 0.000 68.840 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.160 0.000 46.760 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 24.080 0.000 24.680 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 2.000 0.000 2.600 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 49.000 5.000 50.500 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 83.215 189.050 85.225 214.870 ;
        RECT 87.215 189.050 91.175 211.150 ;
        RECT 97.215 189.050 101.175 211.150 ;
        RECT 107.215 189.050 111.175 211.150 ;
        RECT 117.215 189.050 119.225 212.870 ;
      LAYER nwell ;
        RECT 123.215 189.050 127.175 211.240 ;
        RECT 133.215 189.050 137.175 211.240 ;
      LAYER pwell ;
        RECT 141.215 189.050 143.225 212.870 ;
        RECT 149.215 189.050 153.175 211.150 ;
        RECT 160.215 189.050 164.175 211.150 ;
      LAYER nwell ;
        RECT 171.415 200.695 177.775 202.300 ;
      LAYER pwell ;
        RECT 172.550 199.495 176.500 200.175 ;
        RECT 171.755 199.305 171.925 199.475 ;
      LAYER li1 ;
        RECT 83.395 214.520 85.045 214.690 ;
        RECT 83.395 189.400 83.565 214.520 ;
        RECT 84.045 211.880 84.395 214.040 ;
        RECT 84.045 189.880 84.395 192.040 ;
        RECT 84.875 189.400 85.045 214.520 ;
        RECT 117.395 212.520 119.045 212.690 ;
        RECT 83.395 189.230 85.045 189.400 ;
        RECT 87.395 210.800 90.995 210.970 ;
        RECT 87.395 189.400 87.565 210.800 ;
        RECT 88.195 210.290 90.195 210.460 ;
        RECT 87.965 190.080 88.135 210.120 ;
        RECT 90.255 190.080 90.425 210.120 ;
        RECT 88.195 189.740 90.195 189.910 ;
        RECT 90.825 189.400 90.995 210.800 ;
        RECT 87.395 189.230 90.995 189.400 ;
        RECT 97.395 210.800 100.995 210.970 ;
        RECT 97.395 189.400 97.565 210.800 ;
        RECT 98.195 210.290 100.195 210.460 ;
        RECT 97.965 190.080 98.135 210.120 ;
        RECT 100.255 190.080 100.425 210.120 ;
        RECT 98.195 189.740 100.195 189.910 ;
        RECT 100.825 189.400 100.995 210.800 ;
        RECT 97.395 189.230 100.995 189.400 ;
        RECT 107.395 210.800 110.995 210.970 ;
        RECT 107.395 189.400 107.565 210.800 ;
        RECT 108.195 210.290 110.195 210.460 ;
        RECT 107.965 190.080 108.135 210.120 ;
        RECT 110.255 190.080 110.425 210.120 ;
        RECT 108.195 189.740 110.195 189.910 ;
        RECT 110.825 189.400 110.995 210.800 ;
        RECT 107.395 189.230 110.995 189.400 ;
        RECT 117.395 189.400 117.565 212.520 ;
        RECT 118.045 209.880 118.395 212.040 ;
        RECT 118.045 189.880 118.395 192.040 ;
        RECT 118.875 189.400 119.045 212.520 ;
        RECT 141.395 212.520 143.045 212.690 ;
        RECT 117.395 189.230 119.045 189.400 ;
        RECT 123.395 210.890 126.995 211.060 ;
        RECT 123.395 189.400 123.565 210.890 ;
        RECT 124.195 210.380 126.195 210.550 ;
        RECT 123.965 190.125 124.135 210.165 ;
        RECT 126.255 190.125 126.425 210.165 ;
        RECT 126.825 208.420 126.995 210.890 ;
        RECT 133.395 210.890 136.995 211.060 ;
        RECT 133.395 208.420 133.565 210.890 ;
        RECT 134.195 210.380 136.195 210.550 ;
        RECT 126.745 208.080 127.085 208.420 ;
        RECT 133.345 208.080 133.685 208.420 ;
        RECT 124.195 189.740 126.195 189.910 ;
        RECT 126.825 189.400 126.995 208.080 ;
        RECT 123.395 189.230 126.995 189.400 ;
        RECT 133.395 189.400 133.565 208.080 ;
        RECT 133.965 190.125 134.135 210.165 ;
        RECT 136.255 190.125 136.425 210.165 ;
        RECT 134.195 189.740 136.195 189.910 ;
        RECT 136.825 189.400 136.995 210.890 ;
        RECT 133.395 189.230 136.995 189.400 ;
        RECT 141.395 189.400 141.565 212.520 ;
        RECT 142.045 209.880 142.395 212.040 ;
        RECT 142.045 189.880 142.395 192.040 ;
        RECT 142.875 189.400 143.045 212.520 ;
        RECT 141.395 189.230 143.045 189.400 ;
        RECT 149.395 210.800 152.995 210.970 ;
        RECT 149.395 189.400 149.565 210.800 ;
        RECT 150.195 210.290 152.195 210.460 ;
        RECT 149.965 190.080 150.135 210.120 ;
        RECT 152.255 190.080 152.425 210.120 ;
        RECT 150.195 189.740 152.195 189.910 ;
        RECT 152.825 189.400 152.995 210.800 ;
        RECT 149.395 189.230 152.995 189.400 ;
        RECT 160.395 210.800 163.995 210.970 ;
        RECT 160.395 189.400 160.565 210.800 ;
        RECT 161.195 210.290 163.195 210.460 ;
        RECT 160.965 190.080 161.135 210.120 ;
        RECT 163.255 190.080 163.425 210.120 ;
        RECT 161.195 189.740 163.195 189.910 ;
        RECT 163.825 189.400 163.995 210.800 ;
        RECT 171.605 202.025 177.585 202.195 ;
        RECT 171.740 201.190 172.000 202.025 ;
        RECT 172.170 201.020 172.410 201.825 ;
        RECT 172.580 201.190 172.840 202.025 ;
        RECT 173.010 201.020 173.250 201.825 ;
        RECT 173.420 201.190 173.680 202.025 ;
        RECT 173.850 201.020 174.100 201.825 ;
        RECT 174.270 201.190 174.515 202.025 ;
        RECT 174.685 201.020 174.930 201.825 ;
        RECT 175.100 201.190 175.355 202.025 ;
        RECT 175.525 201.020 175.780 201.825 ;
        RECT 175.950 201.190 176.200 202.025 ;
        RECT 176.370 201.020 176.610 201.825 ;
        RECT 176.780 201.190 177.035 202.025 ;
        RECT 171.720 200.950 177.045 201.020 ;
        RECT 171.720 200.850 180.915 200.950 ;
        RECT 171.720 200.255 171.890 200.850 ;
        RECT 172.060 200.425 176.470 200.680 ;
        RECT 176.715 200.255 180.915 200.850 ;
        RECT 171.720 200.150 180.915 200.255 ;
        RECT 171.720 200.085 177.045 200.150 ;
        RECT 172.640 199.475 172.970 199.915 ;
        RECT 173.140 199.670 173.330 200.085 ;
        RECT 173.500 199.475 173.830 199.915 ;
        RECT 174.000 199.670 174.190 200.085 ;
        RECT 174.360 199.475 174.690 199.915 ;
        RECT 174.860 199.670 175.050 200.085 ;
        RECT 175.220 199.475 175.550 199.915 ;
        RECT 175.720 199.670 175.910 200.085 ;
        RECT 176.080 199.475 176.410 199.915 ;
        RECT 171.605 199.305 177.585 199.475 ;
        RECT 160.395 189.230 163.995 189.400 ;
      LAYER mcon ;
        RECT 84.125 211.965 84.315 213.950 ;
        RECT 84.125 189.970 84.315 191.955 ;
        RECT 88.275 210.290 90.115 210.460 ;
        RECT 87.965 190.160 88.135 210.040 ;
        RECT 90.255 190.160 90.425 210.040 ;
        RECT 88.275 189.740 90.115 189.910 ;
        RECT 98.275 210.290 100.115 210.460 ;
        RECT 97.965 190.160 98.135 210.040 ;
        RECT 100.255 190.160 100.425 210.040 ;
        RECT 98.275 189.740 100.115 189.910 ;
        RECT 108.275 210.290 110.115 210.460 ;
        RECT 107.965 190.160 108.135 210.040 ;
        RECT 110.255 190.160 110.425 210.040 ;
        RECT 108.275 189.740 110.115 189.910 ;
        RECT 118.125 209.965 118.315 211.950 ;
        RECT 118.125 189.970 118.315 191.955 ;
        RECT 124.275 210.380 126.115 210.550 ;
        RECT 123.965 190.205 124.135 210.085 ;
        RECT 126.255 190.205 126.425 210.085 ;
        RECT 134.275 210.380 136.115 210.550 ;
        RECT 126.745 208.080 127.085 208.420 ;
        RECT 133.345 208.080 133.685 208.420 ;
        RECT 124.275 189.740 126.115 189.910 ;
        RECT 133.965 190.205 134.135 210.085 ;
        RECT 136.255 190.205 136.425 210.085 ;
        RECT 134.275 189.740 136.115 189.910 ;
        RECT 142.125 209.965 142.315 211.950 ;
        RECT 142.125 189.970 142.315 191.955 ;
        RECT 150.275 210.290 152.115 210.460 ;
        RECT 149.965 190.160 150.135 210.040 ;
        RECT 152.255 190.160 152.425 210.040 ;
        RECT 150.275 189.740 152.115 189.910 ;
        RECT 161.275 210.290 163.115 210.460 ;
        RECT 160.965 190.160 161.135 210.040 ;
        RECT 163.255 190.160 163.425 210.040 ;
        RECT 161.275 189.740 163.115 189.910 ;
        RECT 171.750 202.025 171.920 202.195 ;
        RECT 172.210 202.025 172.380 202.195 ;
        RECT 172.670 202.025 172.840 202.195 ;
        RECT 173.130 202.025 173.300 202.195 ;
        RECT 173.590 202.025 173.760 202.195 ;
        RECT 174.050 202.025 174.220 202.195 ;
        RECT 174.510 202.025 174.680 202.195 ;
        RECT 174.970 202.025 175.140 202.195 ;
        RECT 175.430 202.025 175.600 202.195 ;
        RECT 175.890 202.025 176.060 202.195 ;
        RECT 176.350 202.025 176.520 202.195 ;
        RECT 176.810 202.025 176.980 202.195 ;
        RECT 177.270 202.025 177.440 202.195 ;
        RECT 175.030 200.465 175.200 200.635 ;
        RECT 180.145 200.180 180.885 200.920 ;
        RECT 171.750 199.305 171.920 199.475 ;
        RECT 172.210 199.305 172.380 199.475 ;
        RECT 172.670 199.305 172.840 199.475 ;
        RECT 173.130 199.305 173.300 199.475 ;
        RECT 173.590 199.305 173.760 199.475 ;
        RECT 174.050 199.305 174.220 199.475 ;
        RECT 174.510 199.305 174.680 199.475 ;
        RECT 174.970 199.305 175.140 199.475 ;
        RECT 175.430 199.305 175.600 199.475 ;
        RECT 175.890 199.305 176.060 199.475 ;
        RECT 176.350 199.305 176.520 199.475 ;
        RECT 176.810 199.305 176.980 199.475 ;
        RECT 177.270 199.305 177.440 199.475 ;
      LAYER met1 ;
        RECT 87.115 216.650 171.115 221.050 ;
        RECT 83.715 215.850 171.115 216.650 ;
        RECT 83.720 213.255 84.510 215.850 ;
        RECT 87.115 214.050 171.115 215.850 ;
        RECT 118.015 213.555 118.415 214.050 ;
        RECT 84.095 211.905 84.345 213.255 ;
        RECT 85.415 211.650 99.615 212.450 ;
        RECT 85.415 194.050 86.215 211.650 ;
        RECT 98.915 210.490 99.415 211.650 ;
        RECT 109.065 210.490 109.565 212.330 ;
        RECT 88.215 210.260 90.175 210.490 ;
        RECT 98.215 210.260 100.175 210.490 ;
        RECT 108.215 210.260 110.175 210.490 ;
        RECT 118.015 210.350 118.420 213.555 ;
        RECT 87.935 194.050 88.165 210.100 ;
        RECT 90.225 194.450 90.455 210.100 ;
        RECT 97.935 194.450 98.165 210.100 ;
        RECT 98.915 209.950 99.415 210.260 ;
        RECT 100.225 208.550 100.455 210.100 ;
        RECT 104.325 208.550 104.925 208.580 ;
        RECT 107.935 208.550 108.165 210.100 ;
        RECT 109.065 209.800 109.565 210.260 ;
        RECT 100.115 207.950 108.315 208.550 ;
        RECT 85.415 193.250 88.515 194.050 ;
        RECT 84.095 191.050 84.345 192.015 ;
        RECT 85.415 191.050 86.215 193.250 ;
        RECT 83.915 190.250 86.215 191.050 ;
        RECT 84.095 189.910 84.345 190.250 ;
        RECT 85.415 187.950 86.215 190.250 ;
        RECT 87.935 190.100 88.165 193.250 ;
        RECT 89.515 192.850 98.715 194.450 ;
        RECT 88.715 189.940 89.515 190.250 ;
        RECT 90.225 190.100 90.455 192.850 ;
        RECT 88.215 189.710 90.175 189.940 ;
        RECT 88.715 187.950 89.515 189.710 ;
        RECT 85.415 187.150 89.515 187.950 ;
        RECT 93.515 184.750 95.115 192.850 ;
        RECT 97.935 190.100 98.165 192.850 ;
        RECT 100.225 190.100 100.455 207.950 ;
        RECT 104.325 207.920 104.925 207.950 ;
        RECT 107.935 190.100 108.165 207.950 ;
        RECT 110.225 191.200 110.455 210.100 ;
        RECT 118.095 209.905 118.345 210.350 ;
        RECT 122.515 209.450 122.915 214.050 ;
        RECT 124.215 210.350 126.175 210.580 ;
        RECT 123.935 209.450 124.165 210.145 ;
        RECT 122.515 209.050 124.315 209.450 ;
        RECT 118.095 191.200 118.345 192.015 ;
        RECT 109.965 190.700 118.465 191.200 ;
        RECT 110.225 190.100 110.455 190.700 ;
        RECT 98.215 189.710 100.175 189.940 ;
        RECT 108.215 189.710 110.175 189.940 ;
        RECT 115.865 188.350 116.365 190.700 ;
        RECT 118.095 189.910 118.345 190.700 ;
        RECT 123.935 190.145 124.165 209.050 ;
        RECT 126.225 191.500 126.455 210.145 ;
        RECT 126.715 208.020 127.115 214.050 ;
        RECT 133.315 208.020 133.715 214.050 ;
        RECT 134.215 210.350 136.175 210.580 ;
        RECT 132.035 200.100 132.595 200.600 ;
        RECT 128.165 191.500 128.665 197.930 ;
        RECT 125.965 191.000 128.665 191.500 ;
        RECT 126.225 190.145 126.455 191.000 ;
        RECT 124.965 189.940 125.465 190.100 ;
        RECT 124.215 189.710 126.175 189.940 ;
        RECT 124.965 188.350 125.465 189.710 ;
        RECT 128.165 188.350 128.665 191.000 ;
        RECT 132.065 195.120 132.565 200.100 ;
        RECT 132.065 194.320 132.615 195.120 ;
        RECT 132.065 191.500 132.565 194.320 ;
        RECT 133.935 191.500 134.165 210.145 ;
        RECT 136.225 209.450 136.455 210.145 ;
        RECT 137.715 209.450 138.115 214.050 ;
        RECT 142.015 209.850 142.415 214.050 ;
        RECT 147.415 214.020 147.915 214.050 ;
        RECT 150.935 211.800 151.495 212.300 ;
        RECT 150.965 210.490 151.465 211.800 ;
        RECT 161.965 210.490 162.465 212.180 ;
        RECT 150.215 210.260 152.175 210.490 ;
        RECT 161.215 210.260 163.175 210.490 ;
        RECT 136.115 209.050 138.115 209.450 ;
        RECT 136.225 198.120 136.455 209.050 ;
        RECT 135.815 197.320 137.015 198.120 ;
        RECT 132.065 191.000 134.365 191.500 ;
        RECT 132.065 188.350 132.565 191.000 ;
        RECT 133.935 190.145 134.165 191.000 ;
        RECT 136.225 190.145 136.455 197.320 ;
        RECT 142.095 191.300 142.345 192.015 ;
        RECT 141.965 191.200 144.065 191.300 ;
        RECT 149.935 191.200 150.165 210.100 ;
        RECT 150.965 209.900 151.465 210.260 ;
        RECT 161.965 210.100 162.465 210.260 ;
        RECT 152.225 208.650 152.455 210.100 ;
        RECT 156.285 208.650 156.885 208.680 ;
        RECT 160.935 208.650 161.165 210.100 ;
        RECT 152.015 208.050 161.315 208.650 ;
        RECT 141.965 190.800 150.365 191.200 ;
        RECT 134.215 189.710 136.175 189.940 ;
        RECT 142.095 189.910 142.345 190.800 ;
        RECT 143.565 190.700 150.365 190.800 ;
        RECT 135.065 188.350 135.565 189.710 ;
        RECT 143.565 188.350 144.065 190.700 ;
        RECT 149.935 190.100 150.165 190.700 ;
        RECT 152.225 190.100 152.455 208.050 ;
        RECT 156.285 208.020 156.885 208.050 ;
        RECT 160.935 190.100 161.165 208.050 ;
        RECT 163.225 194.950 163.455 210.100 ;
        RECT 165.415 203.450 167.015 214.050 ;
        RECT 165.315 201.850 179.015 203.450 ;
        RECT 168.815 200.650 169.515 201.050 ;
        RECT 180.815 200.950 186.715 203.050 ;
        RECT 174.970 200.650 175.260 200.665 ;
        RECT 168.815 200.450 175.260 200.650 ;
        RECT 168.815 200.150 169.515 200.450 ;
        RECT 174.970 200.435 175.260 200.450 ;
        RECT 180.085 200.150 186.715 200.950 ;
        RECT 171.605 199.350 177.585 199.630 ;
        RECT 165.215 197.750 178.915 199.350 ;
        RECT 165.215 194.950 166.815 197.750 ;
        RECT 180.815 197.450 186.715 200.150 ;
        RECT 162.515 193.350 166.815 194.950 ;
        RECT 163.225 190.100 163.455 193.350 ;
        RECT 150.215 189.710 152.175 189.940 ;
        RECT 161.215 189.710 163.175 189.940 ;
        RECT 115.865 187.850 128.715 188.350 ;
        RECT 132.015 187.850 144.065 188.350 ;
        RECT 165.215 184.750 166.815 193.350 ;
        RECT 85.615 179.350 169.015 184.750 ;
      LAYER via ;
        RECT 98.915 211.650 99.415 212.150 ;
        RECT 109.065 211.800 109.565 212.300 ;
        RECT 104.325 207.950 104.925 208.550 ;
        RECT 132.065 200.100 132.565 200.600 ;
        RECT 128.165 197.400 128.665 197.900 ;
        RECT 150.965 211.800 151.465 212.300 ;
        RECT 161.965 211.650 162.465 212.150 ;
        RECT 156.285 208.050 156.885 208.650 ;
        RECT 168.865 200.300 169.365 200.800 ;
      LAYER met2 ;
        RECT 146.565 212.800 169.465 213.300 ;
        RECT 146.565 212.300 147.065 212.800 ;
        RECT 150.965 212.300 151.465 212.330 ;
        RECT 98.915 212.150 99.415 212.180 ;
        RECT 98.915 211.650 104.610 212.150 ;
        RECT 109.035 211.800 114.065 212.300 ;
        RECT 98.915 211.620 99.415 211.650 ;
        RECT 104.295 207.950 104.955 208.550 ;
        RECT 104.325 176.180 104.925 207.950 ;
        RECT 113.565 200.600 114.065 211.800 ;
        RECT 146.565 211.800 151.465 212.300 ;
        RECT 155.690 212.150 156.140 212.170 ;
        RECT 132.065 200.600 132.565 200.630 ;
        RECT 113.565 200.100 132.565 200.600 ;
        RECT 132.065 200.070 132.565 200.100 ;
        RECT 146.565 197.900 147.065 211.800 ;
        RECT 150.965 211.770 151.465 211.800 ;
        RECT 155.665 211.650 162.605 212.150 ;
        RECT 155.690 211.630 156.140 211.650 ;
        RECT 168.965 211.140 169.465 212.800 ;
        RECT 168.865 209.800 169.465 211.140 ;
        RECT 156.255 208.050 156.915 208.650 ;
        RECT 128.135 197.400 147.065 197.900 ;
        RECT 104.325 175.580 108.520 176.180 ;
        RECT 156.285 175.200 156.885 208.050 ;
        RECT 168.865 200.270 169.365 209.800 ;
        RECT 156.240 174.600 156.930 175.200 ;
      LAYER via2 ;
        RECT 104.065 211.650 104.565 212.150 ;
        RECT 155.690 211.675 156.140 212.125 ;
        RECT 107.875 175.580 108.475 176.180 ;
        RECT 156.285 174.600 156.885 175.200 ;
      LAYER met3 ;
        RECT 104.040 212.150 104.590 212.175 ;
        RECT 104.040 211.650 156.165 212.150 ;
        RECT 104.040 211.625 104.590 211.650 ;
        RECT 107.850 176.180 108.500 176.205 ;
        RECT 107.850 175.580 110.075 176.180 ;
        RECT 107.850 175.555 108.500 175.580 ;
        RECT 156.260 175.200 156.910 175.225 ;
        RECT 152.225 174.600 156.910 175.200 ;
        RECT 156.260 174.575 156.910 174.600 ;
        RECT 97.615 142.990 129.475 173.390 ;
        RECT 133.995 143.570 165.855 173.970 ;
        RECT 97.615 111.390 129.475 141.790 ;
        RECT 133.995 111.970 165.855 142.370 ;
        RECT 97.615 79.790 129.475 110.190 ;
        RECT 133.995 80.370 165.855 110.770 ;
        RECT 97.615 48.190 129.475 78.590 ;
        RECT 133.995 48.770 165.855 79.170 ;
        RECT 97.615 16.590 129.475 46.990 ;
        RECT 133.995 17.170 165.855 47.570 ;
      LAYER via3 ;
        RECT 109.445 175.580 110.045 176.180 ;
        RECT 152.255 174.600 152.855 175.200 ;
        RECT 129.055 143.130 129.375 173.250 ;
        RECT 165.435 143.710 165.755 173.830 ;
        RECT 129.055 111.530 129.375 141.650 ;
        RECT 165.435 112.110 165.755 142.230 ;
        RECT 129.055 79.930 129.375 110.050 ;
        RECT 165.435 80.510 165.755 110.630 ;
        RECT 129.055 48.330 129.375 78.450 ;
        RECT 165.435 48.910 165.755 79.030 ;
        RECT 129.055 16.730 129.375 46.850 ;
        RECT 165.435 17.310 165.755 47.430 ;
      LAYER met4 ;
        RECT 3.990 223.550 4.290 224.760 ;
        RECT 7.670 223.550 7.970 224.760 ;
        RECT 11.350 223.550 11.650 224.760 ;
        RECT 15.030 223.550 15.330 224.760 ;
        RECT 18.710 223.550 19.010 224.760 ;
        RECT 22.390 223.550 22.690 224.760 ;
        RECT 26.070 223.550 26.370 224.760 ;
        RECT 29.750 223.550 30.050 224.760 ;
        RECT 33.430 223.550 33.730 224.760 ;
        RECT 37.110 223.550 37.410 224.760 ;
        RECT 40.790 223.550 41.090 224.760 ;
        RECT 44.470 223.550 44.770 224.760 ;
        RECT 48.150 223.550 48.450 224.760 ;
        RECT 51.830 223.550 52.130 224.760 ;
        RECT 55.510 223.550 55.810 224.760 ;
        RECT 59.190 223.550 59.490 224.760 ;
        RECT 62.870 223.550 63.170 224.760 ;
        RECT 66.550 223.550 66.850 224.760 ;
        RECT 70.230 223.550 70.530 224.760 ;
        RECT 73.910 223.550 74.210 224.760 ;
        RECT 77.590 223.550 77.890 224.760 ;
        RECT 81.270 223.550 81.570 224.760 ;
        RECT 84.950 223.550 85.250 224.760 ;
        RECT 88.630 223.550 88.930 224.760 ;
        RECT 2.760 222.050 89.560 223.550 ;
        RECT 49.000 220.760 50.500 222.050 ;
        RECT 109.440 176.180 110.050 176.185 ;
        RECT 112.555 176.180 165.865 176.250 ;
        RECT 109.440 175.730 165.865 176.180 ;
        RECT 109.440 175.580 113.385 175.730 ;
        RECT 109.440 175.575 110.050 175.580 ;
        RECT 112.555 172.995 113.075 175.580 ;
        RECT 152.250 175.200 152.860 175.205 ;
        RECT 147.505 175.180 152.860 175.200 ;
        RECT 128.875 174.660 152.860 175.180 ;
        RECT 128.875 173.990 129.395 174.660 ;
        RECT 147.505 174.600 152.860 174.660 ;
        RECT 98.010 143.385 127.620 172.995 ;
        RECT 128.875 168.720 129.475 173.990 ;
        RECT 148.935 173.575 149.455 174.600 ;
        RECT 152.250 174.595 152.860 174.600 ;
        RECT 165.345 174.570 165.865 175.730 ;
        RECT 112.555 141.395 113.075 143.385 ;
        RECT 98.010 111.785 127.620 141.395 ;
        RECT 112.555 109.795 113.075 111.785 ;
        RECT 98.010 80.185 127.620 109.795 ;
        RECT 112.555 78.195 113.075 80.185 ;
        RECT 98.010 48.585 127.620 78.195 ;
        RECT 112.555 46.595 113.075 48.585 ;
        RECT 98.010 16.985 127.620 46.595 ;
        RECT 112.555 15.990 113.075 16.985 ;
        RECT 128.955 15.990 129.475 168.720 ;
        RECT 134.390 143.965 164.000 173.575 ;
        RECT 165.335 168.110 165.865 174.570 ;
        RECT 148.935 141.975 149.455 143.965 ;
        RECT 134.390 112.365 164.000 141.975 ;
        RECT 148.935 110.375 149.455 112.365 ;
        RECT 134.390 80.765 164.000 110.375 ;
        RECT 148.935 78.775 149.455 80.765 ;
        RECT 134.390 49.165 164.000 78.775 ;
        RECT 148.935 47.175 149.455 49.165 ;
        RECT 134.390 17.565 164.000 47.175 ;
        RECT 148.935 16.570 149.455 17.565 ;
        RECT 165.335 16.570 165.855 168.110 ;
  END
END tt_um_mattvenn_relax_osc
END LIBRARY

