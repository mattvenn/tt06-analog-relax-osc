magic
tech sky130A
magscale 1 2
timestamp 1713344109
<< metal1 >>
rect 10916 43408 11216 43414
rect 11216 43108 12388 43408
rect 10916 43102 11216 43108
rect 31312 41214 31432 41748
rect 31306 41094 31312 41214
rect 31432 41094 31438 41214
rect 31044 40438 31050 40498
rect 31110 40438 31116 40498
rect 31050 39646 31110 40438
rect 31312 39204 31432 39210
rect 11556 36112 11856 36118
rect 11856 35812 12520 36112
rect 11556 35806 11856 35812
<< via1 >>
rect 10916 43108 11216 43408
rect 31312 41094 31432 41214
rect 31050 40438 31110 40498
rect 11556 35812 11856 36112
<< metal2 >>
rect 6577 43172 6867 43176
rect 10382 43172 10916 43408
rect 6572 43167 10916 43172
rect 6572 42877 6577 43167
rect 6867 43108 10916 43167
rect 11216 43108 11222 43408
rect 6867 42877 10682 43108
rect 6572 42872 10682 42877
rect 6577 42868 6867 42872
rect 31312 41214 31432 41220
rect 31312 40905 31432 41094
rect 31308 40795 31317 40905
rect 31427 40795 31436 40905
rect 31312 40790 31432 40795
rect 31050 40712 31110 40714
rect 31043 40656 31052 40712
rect 31108 40656 31117 40712
rect 31050 40498 31110 40656
rect 31050 40432 31110 40438
rect 11023 36112 11313 36116
rect 11018 36107 11556 36112
rect 11018 35817 11023 36107
rect 11313 35817 11556 36107
rect 11018 35812 11556 35817
rect 11856 35812 11862 36112
rect 11023 35808 11313 35812
<< via2 >>
rect 6577 42877 6867 43167
rect 31317 40795 31427 40905
rect 31052 40656 31108 40712
rect 11023 35817 11313 36107
<< metal3 >>
rect 5067 43172 5365 43177
rect 5066 43171 6872 43172
rect 5066 42873 5067 43171
rect 5365 43167 6872 43171
rect 5365 42877 6577 43167
rect 6867 42877 6872 43167
rect 5365 42873 6872 42877
rect 5066 42872 6872 42873
rect 5067 42867 5365 42872
rect 31042 40914 31048 40978
rect 31112 40914 31118 40978
rect 31050 40717 31110 40914
rect 31312 40905 31432 40910
rect 31312 40795 31317 40905
rect 31427 40795 31432 40905
rect 31047 40712 31113 40717
rect 31047 40656 31052 40712
rect 31108 40656 31113 40712
rect 31047 40651 31113 40656
rect 31312 40625 31432 40795
rect 31307 40507 31313 40625
rect 31431 40507 31437 40625
rect 31312 40506 31432 40507
rect 10355 36112 10653 36117
rect 10354 36111 11318 36112
rect 10354 35813 10355 36111
rect 10653 36107 11318 36111
rect 10653 35817 11023 36107
rect 11313 35817 11318 36107
rect 10653 35813 11318 35817
rect 10354 35812 11318 35813
rect 10355 35807 10653 35812
<< via3 >>
rect 5067 42873 5365 43171
rect 31048 40914 31112 40978
rect 31313 40507 31431 40625
rect 10355 35813 10653 36111
<< metal4 >>
rect 798 44710 858 45152
rect 1534 44710 1594 45152
rect 2270 44710 2330 45152
rect 3006 44710 3066 45152
rect 3742 44710 3802 45152
rect 4478 44710 4538 45152
rect 5214 44710 5274 45152
rect 5950 44710 6010 45152
rect 6686 44710 6746 45152
rect 7422 44710 7482 45152
rect 8158 44710 8218 45152
rect 8894 44710 8954 45152
rect 9630 44710 9690 45152
rect 10366 44710 10426 45152
rect 11102 44710 11162 45152
rect 11838 44710 11898 45152
rect 12574 44710 12634 45152
rect 13310 44710 13370 45152
rect 14046 44710 14106 45152
rect 14782 44710 14842 45152
rect 15518 44710 15578 45152
rect 16254 44710 16314 45152
rect 16990 44710 17050 45152
rect 552 44410 17484 44710
rect 17726 44612 17786 45152
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 22878 44952 22938 45152
rect 23614 44952 23674 45152
rect 24350 44952 24410 45152
rect 25086 44952 25146 45152
rect 25822 44952 25882 45152
rect 26558 44952 26618 45152
rect 27294 44952 27354 45152
rect 28030 44952 28090 45152
rect 28766 44952 28826 45152
rect 29502 44952 29562 45152
rect 30238 44952 30298 45152
rect 30974 44952 31034 45152
rect 31710 44952 31770 45152
rect 17726 44552 31110 44612
rect 200 43172 500 44152
rect 200 43171 5366 43172
rect 200 42873 5067 43171
rect 5365 42873 5366 43171
rect 200 42872 5366 42873
rect 200 1000 500 42872
rect 9800 36112 10100 44410
rect 31050 40979 31110 44552
rect 31047 40978 31113 40979
rect 31047 40914 31048 40978
rect 31112 40914 31113 40978
rect 31047 40913 31113 40914
rect 31312 40625 31432 40626
rect 31312 40507 31313 40625
rect 31431 40507 31432 40625
rect 9800 36111 10654 36112
rect 9800 35813 10355 36111
rect 10653 35813 10654 36111
rect 9800 35812 10654 35813
rect 9800 1000 10100 35812
rect 400 0 520 200
rect 4816 0 4936 200
rect 9232 0 9352 200
rect 13648 0 13768 200
rect 18064 0 18184 200
rect 22480 0 22600 200
rect 26896 0 27016 200
rect 31312 0 31432 40507
use osc  osc_0 ~/work/asic-workshop/shuttle-2404/tt06-analog-relax-osc/mag
timestamp 1713344109
transform 1 0 7190 0 1 30334
box 3800 -27612 24528 13400
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31312 0 31432 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26896 0 27016 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22480 0 22600 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18064 0 18184 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13648 0 13768 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9232 0 9352 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4816 0 4936 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 400 0 520 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 500 44152 1 FreeSans 2 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 9800 1000 10100 44152 1 FreeSans 2 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
