* NGSPICE file created from osc_parax.ext - technology: sky130A

.subckt osc_parax VSS osc_out osc_a VDD
X0 osc_out.t11 osc_a.t4 VDD.t27 VDD.t26 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X1 osc_out.t12 osc_a.t5 VSS.t17 VSS.t16 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X2 osc_out.t10 osc_a.t6 VDD.t25 VDD.t24 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X3 VDD osc_a VSS.t18 sky130_fd_pr__res_high_po_0p35 l=18
X4 osc_out.t9 osc_a.t7 VDD.t23 VDD.t22 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X5 VDD.t1 osc_b osc_b VDD.t0 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=5.8 ps=40.58 w=20 l=2
**devattr s=232000,8116 d=232000,8116
X6 VDD osc_b VSS.t19 sky130_fd_pr__res_high_po_0p35 l=18
X7 left_cap.t7 right_cap.t6 sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X8 VDD.t21 osc_a.t8 osc_out.t8 VDD.t20 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X9 VSS.t25 cset right_cap.t1 VSS.t24 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=20 l=2
**devattr s=232000,8116 d=232000,8116
X10 left_cap.t7 right_cap.t5 sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X11 VDD.t19 osc_a.t9 osc_out.t7 VDD.t18 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X12 osc_out.t19 osc_a.t10 VSS.t15 VSS.t14 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X13 left_cap.t7 right_cap.t4 sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X14 osc_a.t2 osc_a.t1 VDD.t17 VDD.t16 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=20 l=2
**devattr s=232000,8116 d=232000,8116
X15 VDD.t15 osc_a.t11 osc_out.t6 VDD.t14 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X16 osc_out.t13 osc_a.t12 VSS.t13 VSS.t12 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=4452,274 d=2352,140
X17 right_cap.t7 left_cap.t5 sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X18 osc_a.t0 osc_b left_cap.t0 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=20 l=2
**devattr s=232000,8116 d=232000,8116
X19 VDD cset VSS.t26 sky130_fd_pr__res_high_po_0p35 l=20
X20 VDD.t13 osc_a.t13 osc_out.t5 VDD.t12 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X21 VSS.t11 osc_a.t14 osc_out.t15 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X22 right_cap.t8 left_cap.t6 sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X23 right_cap.t7 left_cap.t4 sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X24 left_cap.t7 right_cap.t3 sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X25 VDD.t7 osc_a.t15 osc_out.t4 VDD.t6 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X26 left_cap.t1 cset VSS.t23 VSS.t22 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=20 l=2
**devattr s=232000,8116 d=232000,8116
X27 VDD.t9 osc_a.t16 osc_out.t3 VDD.t8 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5400,254 d=5500,255
X28 osc_out.t2 osc_a.t17 VDD.t11 VDD.t10 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5500,255 d=5400,254
X29 VSS.t9 osc_a.t18 osc_out.t17 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X30 VSS.t7 osc_a.t19 osc_out.t18 VSS.t6 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=4452,274
X31 right_cap.t7 left_cap.t3 sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X32 VSS.t21 cset cset VSS.t20 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=5.8 ps=40.58 w=20 l=2
**devattr s=232000,8116 d=232000,8116
X33 right_cap.t7 left_cap.t2 sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X34 VSS.t5 osc_a.t20 osc_out.t14 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X35 right_cap.t0 osc_a.t21 osc_b VSS.t3 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=5.8 ps=40.58 w=20 l=2
**devattr s=232000,8116 d=232000,8116
X36 osc_out.t1 osc_a.t22 VDD.t5 VDD.t4 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X37 left_cap.t7 right_cap.t2 sky130_fd_pr__cap_mim_m3_1 l=30 w=30
X38 osc_out.t16 osc_a.t23 VSS.t2 VSS.t1 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
**devattr s=2352,140 d=2352,140
X39 osc_out.t0 osc_a.t24 VDD.t3 VDD.t2 sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
**devattr s=5400,254 d=5400,254
R0 osc_a.n45 osc_a.t21 285.901
R1 osc_a.n48 osc_a.t1 281.341
R2 osc_a.n3 osc_a.t15 225.911
R3 osc_a.n20 osc_a.t4 205.375
R4 osc_a.n4 osc_a.t24 192.8
R5 osc_a.n2 osc_a.t11 192.8
R6 osc_a.n11 osc_a.t6 192.8
R7 osc_a.n14 osc_a.t13 192.8
R8 osc_a.n38 osc_a.t7 192.8
R9 osc_a.n15 osc_a.t8 192.8
R10 osc_a.n31 osc_a.t22 192.8
R11 osc_a.n17 osc_a.t9 192.8
R12 osc_a.n25 osc_a.t17 192.8
R13 osc_a.n19 osc_a.t16 192.8
R14 osc_a.n7 osc_a.n3 169.067
R15 osc_a.n21 osc_a.n20 152
R16 osc_a.n22 osc_a.n18 152
R17 osc_a.n24 osc_a.n23 152
R18 osc_a.n28 osc_a.n27 152
R19 osc_a.n30 osc_a.n29 152
R20 osc_a.n34 osc_a.n33 152
R21 osc_a.n36 osc_a.n35 152
R22 osc_a.n39 osc_a.n1 152
R23 osc_a.n42 osc_a.n41 152
R24 osc_a.n12 osc_a.n0 152
R25 osc_a.n9 osc_a.n8 152
R26 osc_a.n7 osc_a.n6 152
R27 osc_a.n26 osc_a.t12 117.287
R28 osc_a.n16 osc_a.t14 117.287
R29 osc_a.n32 osc_a.t10 117.287
R30 osc_a.n37 osc_a.t18 117.287
R31 osc_a.n40 osc_a.t5 117.287
R32 osc_a.n13 osc_a.t20 117.287
R33 osc_a.n10 osc_a.t23 117.287
R34 osc_a.n5 osc_a.t19 117.287
R35 osc_a.n24 osc_a.n18 28.5014
R36 osc_a.n38 osc_a.n37 24.3101
R37 osc_a.n20 osc_a.n19 22.6335
R38 osc_a.n33 osc_a.n15 21.3762
R39 osc_a.n5 osc_a.n4 20.957
R40 osc_a.n44 osc_a.n43 20.3509
R41 osc_a.n9 osc_a.n2 19.6996
R42 osc_a.n27 osc_a.n26 18.8614
R43 osc_a.n41 osc_a.n40 17.1848
R44 osc_a.n42 osc_a.n1 17.0672
R45 osc_a.n29 osc_a.n28 17.0672
R46 osc_a.n22 osc_a.n21 17.0672
R47 osc_a.n34 osc_a 16.5652
R48 osc_a.n46 osc_a.t2 16.3824
R49 osc_a.n31 osc_a.n30 14.6701
R50 osc_a.n46 osc_a.n45 14.113
R51 osc_a.n8 osc_a 13.5534
R52 osc_a.n11 osc_a.n10 13.4127
R53 osc_a.n48 osc_a.t0 13.3725
R54 osc_a.n12 osc_a.n11 12.9935
R55 osc_a.n14 osc_a.n13 12.5744
R56 osc_a.n35 osc_a 12.5495
R57 osc_a.n23 osc_a 11.5456
R58 osc_a.n23 osc_a 11.5456
R59 osc_a.n40 osc_a.n39 11.317
R60 osc_a.n30 osc_a.n16 11.317
R61 osc_a.n35 osc_a 10.5417
R62 osc_a.n32 osc_a.n31 10.0596
R63 osc_a.n13 osc_a.n12 9.6405
R64 osc_a.n8 osc_a 9.53776
R65 osc_a.n17 osc_a.n16 9.22137
R66 osc_a.n6 osc_a.n2 8.80224
R67 osc_a.n43 osc_a.n0 8.53383
R68 osc_a.n26 osc_a.n25 8.38311
R69 osc_a.n27 osc_a.n17 7.96398
R70 osc_a.n44 osc_a 7.53169
R71 osc_a osc_a.n0 7.52991
R72 osc_a.n36 osc_a.n15 7.12572
R73 osc_a.n43 osc_a 7.02795
R74 osc_a osc_a.n34 6.52599
R75 osc_a.n41 osc_a.n14 6.28746
R76 osc_a.n19 osc_a.n18 5.86833
R77 osc_a.n45 osc_a.n44 5.7255
R78 osc_a.n28 osc_a 5.52207
R79 osc_a osc_a.n22 5.52207
R80 osc_a.n6 osc_a.n5 5.4492
R81 osc_a osc_a.n1 4.51815
R82 osc_a.n37 osc_a.n36 3.77267
R83 osc_a.n33 osc_a.n32 3.77267
R84 osc_a osc_a.n7 3.51423
R85 osc_a.n4 osc_a.n3 2.09615
R86 osc_a.n10 osc_a.n9 2.09615
R87 osc_a osc_a.n42 1.50638
R88 osc_a.n25 osc_a.n24 1.25789
R89 osc_a.n46 osc_a 0.913
R90 osc_a osc_a.n48 0.738
R91 osc_a.n49 osc_a.n47 0.663
R92 osc_a.n29 osc_a 0.502461
R93 osc_a.n21 osc_a 0.502461
R94 osc_a.n39 osc_a.n38 0.41963
R95 osc_a.n47 osc_a 0.146333
R96 osc_a osc_a.n49 0.1255
R97 osc_a.n49 osc_a 0.063
R98 osc_a.n47 osc_a.n46 0.0236481
R99 VDD.n45 VDD.n43 8795.29
R100 VDD.n48 VDD.n47 8795.29
R101 VDD.n37 VDD.n36 8795.29
R102 VDD.n34 VDD.n32 8795.29
R103 VDD.n44 VDD.n40 938.165
R104 VDD.n44 VDD.n41 938.165
R105 VDD.n49 VDD.n41 938.165
R106 VDD.n33 VDD.n29 938.165
R107 VDD.n33 VDD.n30 938.165
R108 VDD.n38 VDD.n30 938.165
R109 VDD.n50 VDD.n49 603.86
R110 VDD.n39 VDD.n38 603.86
R111 VDD.n27 VDD 438.041
R112 VDD.n11 VDD.t7 349.707
R113 VDD.n26 VDD.t27 343.652
R114 VDD.n50 VDD.n40 321.507
R115 VDD.n39 VDD.n29 321.507
R116 VDD.n6 VDD.n5 318.558
R117 VDD.n10 VDD.n9 318.038
R118 VDD.n14 VDD.n8 317.538
R119 VDD.n2 VDD.n1 317.058
R120 VDD.n20 VDD.n4 317.058
R121 VDD.t8 VDD.t10 251.559
R122 VDD.t2 VDD.t6 248.599
R123 VDD.t14 VDD.t2 248.599
R124 VDD.t24 VDD.t14 248.599
R125 VDD.t12 VDD.t24 248.599
R126 VDD.t22 VDD.t12 248.599
R127 VDD.t20 VDD.t22 248.599
R128 VDD.t4 VDD.t20 248.599
R129 VDD.t18 VDD.t4 248.599
R130 VDD.t10 VDD.t18 248.599
R131 VDD.t26 VDD.t8 248.599
R132 VDD VDD.t26 189.409
R133 VDD.n46 VDD.n45 75.6006
R134 VDD.n48 VDD.n42 75.6006
R135 VDD.n37 VDD.n31 75.6006
R136 VDD.n35 VDD.n34 75.6006
R137 VDD.n16 VDD.n15 34.6358
R138 VDD.n20 VDD.n19 34.2593
R139 VDD.n13 VDD.n10 32.7534
R140 VDD.n21 VDD.n2 28.2358
R141 VDD.n1 VDD.t9 27.5805
R142 VDD.n1 VDD.t11 26.5955
R143 VDD.n4 VDD.t5 26.5955
R144 VDD.n4 VDD.t19 26.5955
R145 VDD.n5 VDD.t23 26.5955
R146 VDD.n5 VDD.t21 26.5955
R147 VDD.n8 VDD.t25 26.5955
R148 VDD.n8 VDD.t13 26.5955
R149 VDD.n9 VDD.t3 26.5955
R150 VDD.n9 VDD.t15 26.5955
R151 VDD.n43 VDD.n40 23.1255
R152 VDD.n47 VDD.n41 23.1255
R153 VDD.n32 VDD.n29 23.1255
R154 VDD.n36 VDD.n30 23.1255
R155 VDD.n43 VDD.n42 22.8671
R156 VDD.n47 VDD.n46 22.8671
R157 VDD.n32 VDD.n31 22.8671
R158 VDD.n36 VDD.n35 22.8671
R159 VDD.n26 VDD.n25 22.2123
R160 VDD.n25 VDD.n2 21.4593
R161 VDD.n54 VDD.t1 18.4534
R162 VDD.n51 VDD.t17 18.3784
R163 VDD.n27 VDD.n26 16.5652
R164 VDD.n21 VDD.n20 15.4358
R165 VDD.n14 VDD.n13 12.0476
R166 VDD.n52 VDD.n50 11.113
R167 VDD.n53 VDD.n39 11.113
R168 VDD.n19 VDD.n6 10.1652
R169 VDD.n13 VDD.n12 9.3005
R170 VDD.n15 VDD.n7 9.3005
R171 VDD.n17 VDD.n16 9.3005
R172 VDD.n19 VDD.n18 9.3005
R173 VDD.n20 VDD.n3 9.3005
R174 VDD.n22 VDD.n21 9.3005
R175 VDD.n23 VDD.n2 9.3005
R176 VDD.n25 VDD.n24 9.3005
R177 VDD.n26 VDD.n0 9.3005
R178 VDD.n28 VDD.n27 9.3005
R179 VDD.n11 VDD.n10 6.33664
R180 VDD.n16 VDD.n6 6.02403
R181 VDD.n15 VDD.n14 3.38874
R182 VDD.n45 VDD.n44 3.03329
R183 VDD.n49 VDD.n48 3.03329
R184 VDD.n34 VDD.n33 3.03329
R185 VDD.n38 VDD.n37 3.03329
R186 VDD VDD.n54 1.71914
R187 VDD.n51 VDD 0.586214
R188 VDD.n12 VDD.n11 0.479734
R189 VDD.t16 VDD.n42 0.19977
R190 VDD.n46 VDD.t16 0.19977
R191 VDD.n35 VDD.t0 0.19977
R192 VDD.t0 VDD.n31 0.19977
R193 VDD.n53 VDD.n52 0.118357
R194 VDD.n54 VDD.n53 0.0790714
R195 VDD.n52 VDD.n51 0.0755
R196 VDD.n12 VDD.n7 0.0364375
R197 VDD.n17 VDD.n7 0.0364375
R198 VDD.n18 VDD.n17 0.0364375
R199 VDD.n18 VDD.n3 0.0364375
R200 VDD.n22 VDD.n3 0.0364375
R201 VDD.n23 VDD.n22 0.0364375
R202 VDD.n24 VDD.n23 0.0364375
R203 VDD.n24 VDD.n0 0.0364375
R204 VDD.n28 VDD 0.0184687
R205 VDD VDD.n28 0.009875
R206 VDD.n0 VDD 0.00675
R207 osc_out.n9 osc_out.n8 317.498
R208 osc_out.n11 osc_out.n10 313.452
R209 osc_out.n19 osc_out.n18 313.452
R210 osc_out.n15 osc_out.n14 313.026
R211 osc_out.n13 osc_out.n12 312.618
R212 osc_out.n17 osc_out.n16 312.226
R213 osc_out.n1 osc_out.n0 207.569
R214 osc_out.n3 osc_out.n2 207.569
R215 osc_out.n5 osc_out.n4 207.569
R216 osc_out.n7 osc_out.n6 207.569
R217 osc_out.n9 osc_out.n7 172.8
R218 osc_out.n21 osc_out.n1 60.6123
R219 osc_out.n20 osc_out 57.8991
R220 osc_out.n3 osc_out.n1 50.4476
R221 osc_out.n5 osc_out.n3 50.4476
R222 osc_out.n7 osc_out.n5 50.4476
R223 osc_out.n11 osc_out.n9 45.177
R224 osc_out.n13 osc_out.n11 45.177
R225 osc_out.n17 osc_out.n15 44.8005
R226 osc_out.n19 osc_out.n17 44.424
R227 osc_out.n15 osc_out.n13 44.0476
R228 osc_out.n0 osc_out.t18 40.0005
R229 osc_out.n0 osc_out.t16 40.0005
R230 osc_out.n2 osc_out.t14 40.0005
R231 osc_out.n2 osc_out.t12 40.0005
R232 osc_out.n4 osc_out.t17 40.0005
R233 osc_out.n4 osc_out.t19 40.0005
R234 osc_out.n6 osc_out.t15 40.0005
R235 osc_out.n6 osc_out.t13 40.0005
R236 osc_out.n8 osc_out.t3 26.5955
R237 osc_out.n8 osc_out.t11 26.5955
R238 osc_out.n10 osc_out.t7 26.5955
R239 osc_out.n10 osc_out.t2 26.5955
R240 osc_out.n12 osc_out.t8 26.5955
R241 osc_out.n12 osc_out.t1 26.5955
R242 osc_out.n14 osc_out.t5 26.5955
R243 osc_out.n14 osc_out.t9 26.5955
R244 osc_out.n16 osc_out.t6 26.5955
R245 osc_out.n16 osc_out.t10 26.5955
R246 osc_out.n18 osc_out.t4 26.5955
R247 osc_out.n18 osc_out.t0 26.5955
R248 osc_out.n21 osc_out 12.6066
R249 osc_out osc_out.n19 11.7852
R250 osc_out.n20 osc_out 11.055
R251 osc_out osc_out.n20 2.13383
R252 osc_out osc_out.n21 0.582318
R253 VSS.n83 VSS.n31 16164.9
R254 VSS.n52 VSS.n44 15412.4
R255 VSS.n48 VSS.n44 15412.4
R256 VSS.n52 VSS.n45 15412.4
R257 VSS.n59 VSS.n41 14386.8
R258 VSS.n55 VSS.n41 14386.8
R259 VSS.n59 VSS.n42 14386.8
R260 VSS.n55 VSS.n42 14386.8
R261 VSS.n66 VSS.n38 14386.8
R262 VSS.n62 VSS.n38 14386.8
R263 VSS.n66 VSS.n39 14386.8
R264 VSS.n62 VSS.n39 14386.8
R265 VSS.n74 VSS.n35 14386.8
R266 VSS.n70 VSS.n35 14386.8
R267 VSS.n74 VSS.n36 14386.8
R268 VSS.n70 VSS.n36 14386.8
R269 VSS.n96 VSS.n91 14386.8
R270 VSS.n91 VSS.n27 14386.8
R271 VSS.n27 VSS.n25 14386.8
R272 VSS.n96 VSS.n25 14386.8
R273 VSS.n100 VSS.n21 14386.8
R274 VSS.n100 VSS.n22 14386.8
R275 VSS.n104 VSS.n22 14386.8
R276 VSS.n104 VSS.n21 14386.8
R277 VSS.n81 VSS.n32 14253.5
R278 VSS.n77 VSS.n32 14253.5
R279 VSS.n81 VSS.n33 14253.5
R280 VSS.n77 VSS.n33 14253.5
R281 VSS.n89 VSS.n28 14253.5
R282 VSS.n85 VSS.n28 14253.5
R283 VSS.n89 VSS.n29 14253.5
R284 VSS.n85 VSS.n29 14253.5
R285 VSS.t24 VSS.t6 7711.91
R286 VSS.n84 VSS.n83 4061.27
R287 VSS.n83 VSS.n82 3715.75
R288 VSS.n106 VSS.n105 2820.61
R289 VSS.t19 VSS.n26 2743.15
R290 VSS.n99 VSS.n98 2423.87
R291 VSS.t3 VSS.n90 1780.1
R292 VSS.n98 VSS.t24 1757.41
R293 VSS.n107 VSS.n106 1198.25
R294 VSS.n51 VSS.n46 1001.41
R295 VSS.n49 VSS.n46 1001.41
R296 VSS.n51 VSS.n50 1001.41
R297 VSS.n50 VSS.n49 1001.41
R298 VSS.n58 VSS.n43 934.777
R299 VSS.n56 VSS.n43 934.777
R300 VSS.n58 VSS.n57 934.777
R301 VSS.n57 VSS.n56 934.777
R302 VSS.n65 VSS.n40 934.777
R303 VSS.n63 VSS.n40 934.777
R304 VSS.n65 VSS.n64 934.777
R305 VSS.n64 VSS.n63 934.777
R306 VSS.n73 VSS.n37 934.777
R307 VSS.n71 VSS.n37 934.777
R308 VSS.n73 VSS.n72 934.777
R309 VSS.n72 VSS.n71 934.777
R310 VSS.n95 VSS.n94 934.777
R311 VSS.n94 VSS.n93 934.777
R312 VSS.n93 VSS.n92 934.777
R313 VSS.n95 VSS.n92 934.777
R314 VSS.n101 VSS.n23 934.777
R315 VSS.n102 VSS.n101 934.777
R316 VSS.n103 VSS.n102 934.777
R317 VSS.n103 VSS.n23 934.777
R318 VSS.n80 VSS.n34 926.119
R319 VSS.n78 VSS.n34 926.119
R320 VSS.n80 VSS.n79 926.119
R321 VSS.n79 VSS.n78 926.119
R322 VSS.n88 VSS.n30 926.119
R323 VSS.n86 VSS.n30 926.119
R324 VSS.n88 VSS.n87 926.119
R325 VSS.n87 VSS.n86 926.119
R326 VSS.n76 VSS.n75 903.375
R327 VSS.n61 VSS.n60 903.375
R328 VSS.n31 VSS.n24 809.014
R329 VSS.n68 VSS.n31 685.96
R330 VSS.n105 VSS.t24 648.004
R331 VSS.t3 VSS.n26 648.004
R332 VSS.n69 VSS.n68 586.438
R333 VSS.n99 VSS.n24 579.991
R334 VSS.t12 VSS 477.974
R335 VSS.n54 VSS.n53 346.5
R336 VSS.n68 VSS.n67 316.938
R337 VSS.n30 VSS.n28 292.5
R338 VSS.n28 VSS.t19 292.5
R339 VSS.n79 VSS.n33 292.5
R340 VSS.n33 VSS.t18 292.5
R341 VSS.n34 VSS.n32 292.5
R342 VSS.n32 VSS.t18 292.5
R343 VSS.n50 VSS.n45 292.5
R344 VSS.n46 VSS.n44 292.5
R345 VSS.n44 VSS.t26 292.5
R346 VSS.n87 VSS.n29 292.5
R347 VSS.n29 VSS.t19 292.5
R348 VSS.n47 VSS.n45 285.058
R349 VSS.n5 VSS.t7 245.403
R350 VSS.n16 VSS.t13 240.127
R351 VSS.n97 VSS.t3 235.814
R352 VSS.n75 VSS.t0 235.812
R353 VSS.n69 VSS.t0 235.812
R354 VSS.n67 VSS.t22 235.812
R355 VSS.n61 VSS.t22 235.812
R356 VSS.n60 VSS.t20 235.812
R357 VSS.n54 VSS.t20 235.812
R358 VSS.n7 VSS.n6 200.127
R359 VSS.n10 VSS.n9 200.127
R360 VSS.n14 VSS.n3 200.127
R361 VSS.n97 VSS.n25 175.472
R362 VSS.t6 VSS.t1 162.474
R363 VSS.t1 VSS.t4 162.474
R364 VSS.t4 VSS.t16 162.474
R365 VSS.t16 VSS.t8 162.474
R366 VSS.t8 VSS.t14 162.474
R367 VSS.t14 VSS.t10 162.474
R368 VSS.t10 VSS.t12 162.474
R369 VSS.n90 VSS.t19 159.962
R370 VSS.n84 VSS.t19 159.962
R371 VSS.n98 VSS.n97 158.814
R372 VSS.n106 VSS 143.582
R373 VSS.n48 VSS.n47 107.081
R374 VSS.n82 VSS.t18 101.751
R375 VSS.n76 VSS.t18 101.751
R376 VSS.n53 VSS.t26 101.751
R377 VSS.n23 VSS.n21 73.1255
R378 VSS.n21 VSS.t24 73.1255
R379 VSS.n96 VSS.n95 73.1255
R380 VSS.t3 VSS.n96 73.1255
R381 VSS.n72 VSS.n36 73.1255
R382 VSS.n36 VSS.t0 73.1255
R383 VSS.n37 VSS.n35 73.1255
R384 VSS.n35 VSS.t0 73.1255
R385 VSS.n64 VSS.n39 73.1255
R386 VSS.n39 VSS.t22 73.1255
R387 VSS.n40 VSS.n38 73.1255
R388 VSS.n38 VSS.t22 73.1255
R389 VSS.n57 VSS.n42 73.1255
R390 VSS.n42 VSS.t20 73.1255
R391 VSS.n43 VSS.n41 73.1255
R392 VSS.n41 VSS.t20 73.1255
R393 VSS.n102 VSS.n22 73.1255
R394 VSS.n22 VSS.t24 73.1255
R395 VSS.n93 VSS.n27 73.1255
R396 VSS.t3 VSS.n27 73.1255
R397 VSS.n24 VSS.t24 68.0125
R398 VSS.n6 VSS.t2 40.0005
R399 VSS.n6 VSS.t5 40.0005
R400 VSS.n9 VSS.t17 40.0005
R401 VSS.n9 VSS.t9 40.0005
R402 VSS.n3 VSS.t15 40.0005
R403 VSS.n3 VSS.t11 40.0005
R404 VSS.n20 VSS.n0 34.6358
R405 VSS.n10 VSS.n8 27.4829
R406 VSS.n16 VSS.n0 25.977
R407 VSS.n107 VSS.n20 23.7181
R408 VSS.n14 VSS.n2 22.9652
R409 VSS.n15 VSS.n14 21.4593
R410 VSS.n16 VSS.n15 18.4476
R411 VSS.n10 VSS.n2 16.9417
R412 VSS.n8 VSS.n7 12.424
R413 VSS.n71 VSS.n70 9.59066
R414 VSS.n70 VSS.n69 9.59066
R415 VSS.n74 VSS.n73 9.59066
R416 VSS.n75 VSS.n74 9.59066
R417 VSS.n63 VSS.n62 9.59066
R418 VSS.n62 VSS.n61 9.59066
R419 VSS.n66 VSS.n65 9.59066
R420 VSS.n67 VSS.n66 9.59066
R421 VSS.n56 VSS.n55 9.59066
R422 VSS.n55 VSS.n54 9.59066
R423 VSS.n59 VSS.n58 9.59066
R424 VSS.n60 VSS.n59 9.59066
R425 VSS.n101 VSS.n100 9.59066
R426 VSS.n100 VSS.n99 9.59066
R427 VSS.n104 VSS.n103 9.59066
R428 VSS.n105 VSS.n104 9.59066
R429 VSS.n94 VSS.n91 9.59066
R430 VSS.n91 VSS.n26 9.59066
R431 VSS.n92 VSS.n25 9.59066
R432 VSS.n108 VSS.n107 9.3005
R433 VSS.n8 VSS.n4 9.3005
R434 VSS.n11 VSS.n10 9.3005
R435 VSS.n12 VSS.n2 9.3005
R436 VSS.n14 VSS.n13 9.3005
R437 VSS.n15 VSS.n1 9.3005
R438 VSS.n17 VSS.n16 9.3005
R439 VSS.n18 VSS.n0 9.3005
R440 VSS.n20 VSS.n19 9.3005
R441 VSS.n86 VSS.n85 8.86414
R442 VSS.n85 VSS.n84 8.86414
R443 VSS.n89 VSS.n88 8.86414
R444 VSS.n90 VSS.n89 8.86414
R445 VSS.n78 VSS.n77 8.86414
R446 VSS.n77 VSS.n76 8.86414
R447 VSS.n81 VSS.n80 8.86414
R448 VSS.n82 VSS.n81 8.86414
R449 VSS.n49 VSS.n48 8.1255
R450 VSS.n52 VSS.n51 8.1255
R451 VSS.n53 VSS.n52 8.1255
R452 VSS.n109 VSS.t21 7.61045
R453 VSS.n109 VSS.t23 7.5917
R454 VSS.n111 VSS.t25 7.23714
R455 VSS.n7 VSS.n5 6.81933
R456 VSS.n111 VSS.n110 2.3321
R457 VSS.n47 VSS.t26 2.03318
R458 VSS.n5 VSS.n4 0.688483
R459 VSS.n110 VSS.n109 0.633312
R460 VSS VSS.n111 0.620031
R461 VSS.n110 VSS 0.157907
R462 VSS.n11 VSS.n4 0.0310851
R463 VSS.n12 VSS.n11 0.0310851
R464 VSS.n13 VSS.n12 0.0310851
R465 VSS.n13 VSS.n1 0.0310851
R466 VSS.n17 VSS.n1 0.0310851
R467 VSS.n18 VSS.n17 0.0310851
R468 VSS.n19 VSS.n18 0.0310851
R469 VSS.n108 VSS 0.0157926
R470 VSS VSS.n108 0.00881117
R471 VSS.n19 VSS 0.00581915
R472 left_cap.n1 left_cap.t1 9.38826
R473 left_cap.n1 left_cap.t0 9.20909
R474 left_cap left_cap.n0 7.91907
R475 left_cap left_cap.n1 7.80107
R476 left_cap.n0 left_cap.t6 6.28228
R477 left_cap.t5 left_cap.t3 2.92748
R478 left_cap.t6 left_cap.t2 2.85665
R479 left_cap.t2 left_cap.t4 2.85665
R480 left_cap.t4 left_cap.t5 2.85665
R481 left_cap.n0 left_cap.t7 0.93824
R482 right_cap.n0 right_cap.t1 9.48011
R483 right_cap.n0 right_cap.t0 9.43427
R484 right_cap right_cap.n0 8.02607
R485 right_cap right_cap.t8 7.45138
R486 right_cap.t8 right_cap.t2 3.21837
R487 right_cap.t6 right_cap.t3 2.92748
R488 right_cap.t2 right_cap.t5 2.85665
R489 right_cap.t5 right_cap.t4 2.85665
R490 right_cap.t4 right_cap.t6 2.85665
R491 right_cap.t8 right_cap.t7 1.02493
C0 left_cap cset 0.733616f
C1 right_cap cset 0.732846f
C2 osc_a left_cap 0.615488f
C3 osc_a right_cap 0.732557f
C4 left_cap osc_b 0.74314f
C5 osc_b right_cap 0.616311f
C6 left_cap right_cap 0.798551p
C7 VDD osc_out 1.21047f
C8 VDD cset 1.83901f
C9 osc_a VDD 6.22817f
C10 osc_a osc_out 1.44545f
C11 osc_a cset 1.10628f
C12 VDD osc_b 4.08243f
C13 osc_b cset 0.550344f
C14 VDD left_cap 0.063197f
C15 osc_a osc_b 2.2743f
C16 VDD right_cap 0.07197f
C17 osc_out VSS 2.85407f
C18 osc_a VSS 18.50762f
C19 VDD VSS 58.746506f
C20 right_cap VSS 93.06754f
C21 osc_b VSS 10.9295f
C22 left_cap VSS 0.101902p
C23 cset VSS 17.3869f
C24 right_cap.t7 VSS 0.284166p
C25 right_cap.t8 VSS 0.227929p
C26 right_cap.t3 VSS 56.5149f
C27 right_cap.t6 VSS 56.817f
C28 right_cap.t4 VSS 56.666f
C29 right_cap.t5 VSS 56.666f
C30 right_cap.t2 VSS 56.7594f
C31 right_cap.t1 VSS 0.536933f
C32 right_cap.t0 VSS 0.535327f
C33 right_cap.n0 VSS 1.2457f
C34 left_cap.t7 VSS 0.362111p
C35 left_cap.n0 VSS 0.149859p
C36 left_cap.t3 VSS 56.4468f
C37 left_cap.t5 VSS 56.7485f
C38 left_cap.t4 VSS 56.5977f
C39 left_cap.t2 VSS 56.5977f
C40 left_cap.t6 VSS 57.1758f
C41 left_cap.t0 VSS 0.526352f
C42 left_cap.t1 VSS 0.533095f
C43 left_cap.n1 VSS 1.19422f
C44 VDD.t6 VSS 0.023731f
C45 VDD.t2 VSS 0.007756f
C46 VDD.t14 VSS 0.007756f
C47 VDD.t24 VSS 0.007756f
C48 VDD.t12 VSS 0.007756f
C49 VDD.t22 VSS 0.007756f
C50 VDD.t20 VSS 0.007756f
C51 VDD.t4 VSS 0.007756f
C52 VDD.t18 VSS 0.007756f
C53 VDD.t10 VSS 0.007802f
C54 VDD.t8 VSS 0.007802f
C55 VDD.t26 VSS 0.006833f
C56 VDD.n0 VSS 0.004971f
C57 VDD.t27 VSS 0.002971f
C58 VDD.t11 VSS 7.77e-19
C59 VDD.t9 VSS 8.05e-19
C60 VDD.n1 VSS 0.001746f
C61 VDD.n2 VSS 0.003489f
C62 VDD.n3 VSS 0.008469f
C63 VDD.t5 VSS 7.77e-19
C64 VDD.t19 VSS 7.77e-19
C65 VDD.n4 VSS 0.001717f
C66 VDD.t23 VSS 7.77e-19
C67 VDD.t21 VSS 7.77e-19
C68 VDD.n5 VSS 0.001716f
C69 VDD.n6 VSS 0.00288f
C70 VDD.n7 VSS 0.008469f
C71 VDD.t25 VSS 7.77e-19
C72 VDD.t13 VSS 7.77e-19
C73 VDD.n8 VSS 0.001717f
C74 VDD.t3 VSS 7.77e-19
C75 VDD.t15 VSS 7.77e-19
C76 VDD.n9 VSS 0.001716f
C77 VDD.n10 VSS 0.003521f
C78 VDD.t7 VSS 0.003041f
C79 VDD.n11 VSS 0.01004f
C80 VDD.n12 VSS 0.06337f
C81 VDD.n13 VSS 5.82e-19
C82 VDD.n14 VSS 0.002986f
C83 VDD.n15 VSS 4.94e-19
C84 VDD.n16 VSS 5.28e-19
C85 VDD.n17 VSS 0.008469f
C86 VDD.n18 VSS 0.008469f
C87 VDD.n19 VSS 5.77e-19
C88 VDD.n20 VSS 0.003489f
C89 VDD.n21 VSS 5.67e-19
C90 VDD.n22 VSS 0.008469f
C91 VDD.n23 VSS 0.008469f
C92 VDD.n24 VSS 0.008469f
C93 VDD.n25 VSS 5.67e-19
C94 VDD.n26 VSS 0.003531f
C95 VDD.n27 VSS 0.011317f
C96 VDD.n28 VSS 0.003222f
C97 VDD.t1 VSS 0.083682f
C98 VDD.n29 VSS 0.01661f
C99 VDD.n30 VSS 0.024659f
C100 VDD.n32 VSS 0.024659f
C101 VDD.n33 VSS 0.024418f
C102 VDD.n34 VSS 0.299648f
C103 VDD.t0 VSS 0.460613f
C104 VDD.n36 VSS 0.024659f
C105 VDD.n37 VSS 0.299648f
C106 VDD.n38 VSS 0.020055f
C107 VDD.n39 VSS 0.015426f
C108 VDD.n40 VSS 0.01661f
C109 VDD.n41 VSS 0.024659f
C110 VDD.n43 VSS 0.024659f
C111 VDD.n44 VSS 0.024418f
C112 VDD.n45 VSS 0.299648f
C113 VDD.t16 VSS 0.460613f
C114 VDD.n47 VSS 0.024659f
C115 VDD.n48 VSS 0.299648f
C116 VDD.n49 VSS 0.020055f
C117 VDD.n50 VSS 0.015426f
C118 VDD.t17 VSS 0.093994f
C119 VDD.n51 VSS 1.59338f
C120 VDD.n52 VSS 0.460335f
C121 VDD.n53 VSS 0.46839f
C122 VDD.n54 VSS 2.59477f
C123 osc_a.n0 VSS 0.001627f
C124 osc_a.n1 VSS 0.002186f
C125 osc_a.t13 VSS 0.004007f
C126 osc_a.t20 VSS 0.00157f
C127 osc_a.t6 VSS 0.004007f
C128 osc_a.t23 VSS 0.00157f
C129 osc_a.t11 VSS 0.004007f
C130 osc_a.n2 VSS 0.005691f
C131 osc_a.t15 VSS 0.005186f
C132 osc_a.n3 VSS 0.01202f
C133 osc_a.t19 VSS 0.00157f
C134 osc_a.t24 VSS 0.004007f
C135 osc_a.n4 VSS 0.004946f
C136 osc_a.n5 VSS 0.004702f
C137 osc_a.n6 VSS 0.001948f
C138 osc_a.n7 VSS 0.005147f
C139 osc_a.n8 VSS 0.002339f
C140 osc_a.n9 VSS 0.002979f
C141 osc_a.n10 VSS 0.003212f
C142 osc_a.n11 VSS 0.005405f
C143 osc_a.n12 VSS 0.003094f
C144 osc_a.n13 VSS 0.004129f
C145 osc_a.n14 VSS 0.004373f
C146 osc_a.t5 VSS 0.00157f
C147 osc_a.t7 VSS 0.004007f
C148 osc_a.t18 VSS 0.00157f
C149 osc_a.t8 VSS 0.004007f
C150 osc_a.n15 VSS 0.005691f
C151 osc_a.t10 VSS 0.00157f
C152 osc_a.t22 VSS 0.004007f
C153 osc_a.t14 VSS 0.00157f
C154 osc_a.n16 VSS 0.0039f
C155 osc_a.t9 VSS 0.004007f
C156 osc_a.n17 VSS 0.004144f
C157 osc_a.t12 VSS 0.00157f
C158 osc_a.t17 VSS 0.004007f
C159 osc_a.n18 VSS 0.0047f
C160 osc_a.t16 VSS 0.004007f
C161 osc_a.n19 VSS 0.005692f
C162 osc_a.t4 VSS 0.004328f
C163 osc_a.n20 VSS 0.009727f
C164 osc_a.n21 VSS 0.001779f
C165 osc_a.n22 VSS 0.002288f
C166 osc_a.n23 VSS 0.002339f
C167 osc_a.n24 VSS 0.004069f
C168 osc_a.n25 VSS 0.003112f
C169 osc_a.n26 VSS 0.004817f
C170 osc_a.n27 VSS 0.003667f
C171 osc_a.n28 VSS 0.002288f
C172 osc_a.n29 VSS 0.001779f
C173 osc_a.n30 VSS 0.003553f
C174 osc_a.n31 VSS 0.005175f
C175 osc_a.n32 VSS 0.002982f
C176 osc_a.n33 VSS 0.003438f
C177 osc_a.n34 VSS 0.002339f
C178 osc_a.n35 VSS 0.002339f
C179 osc_a.n36 VSS 0.001489f
C180 osc_a.n37 VSS 0.004931f
C181 osc_a.n38 VSS 0.005175f
C182 osc_a.n39 VSS 0.001604f
C183 osc_a.n40 VSS 0.004988f
C184 osc_a.n41 VSS 0.003209f
C185 osc_a.n42 VSS 0.001881f
C186 osc_a.n43 VSS 0.050916f
C187 osc_a.n44 VSS 0.659076f
C188 osc_a.t21 VSS 1.29569f
C189 osc_a.n45 VSS 1.21696f
C190 osc_a.t2 VSS 0.29417f
C191 osc_a.n46 VSS 0.616766f
C192 osc_a.n47 VSS 0.215047f
C193 osc_a.t1 VSS 1.29256f
C194 osc_a.t0 VSS 0.481708f
C195 osc_a.n48 VSS 0.879669f
C196 osc_a.n49 VSS 0.039873f
.ends

