VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO osc
  CLASS BLOCK ;
  FOREIGN osc ;
  ORIGIN -19.000 138.060 ;
  SIZE 103.500 BY 205.060 ;
  PIN osc_out
    ANTENNADIFFAREA 2.090400 ;
    PORT
      LAYER met1 ;
        RECT 116.900 46.200 117.900 47.200 ;
    END
  END osc_out
  PIN VDD
    ANTENNADIFFAREA 30.536200 ;
    PORT
      LAYER met1 ;
        RECT 25.700 62.500 26.700 63.500 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 17.975399 ;
    PORT
      LAYER met1 ;
        RECT 23.300 26.800 24.300 27.800 ;
    END
  END VSS
  OBS
      LAYER pwell ;
        RECT 19.000 35.000 21.010 60.820 ;
        RECT 23.000 35.000 26.960 57.100 ;
        RECT 33.000 35.000 36.960 57.100 ;
        RECT 43.000 35.000 46.960 57.100 ;
        RECT 53.000 35.000 55.010 58.820 ;
      LAYER nwell ;
        RECT 59.000 35.000 62.960 57.190 ;
        RECT 69.000 35.000 72.960 57.190 ;
      LAYER pwell ;
        RECT 77.000 35.000 79.010 58.820 ;
        RECT 85.000 35.000 88.960 57.100 ;
        RECT 96.000 35.000 99.960 57.100 ;
      LAYER nwell ;
        RECT 107.200 46.645 113.560 48.250 ;
      LAYER pwell ;
        RECT 108.335 45.445 112.285 46.125 ;
        RECT 107.540 45.255 107.710 45.425 ;
      LAYER li1 ;
        RECT 19.180 60.470 20.830 60.640 ;
        RECT 19.180 35.350 19.350 60.470 ;
        RECT 19.830 57.830 20.180 59.990 ;
        RECT 19.830 35.830 20.180 37.990 ;
        RECT 20.660 35.350 20.830 60.470 ;
        RECT 53.180 58.470 54.830 58.640 ;
        RECT 19.180 35.180 20.830 35.350 ;
        RECT 23.180 56.750 26.780 56.920 ;
        RECT 23.180 35.350 23.350 56.750 ;
        RECT 23.980 56.240 25.980 56.410 ;
        RECT 23.750 36.030 23.920 56.070 ;
        RECT 26.040 36.030 26.210 56.070 ;
        RECT 23.980 35.690 25.980 35.860 ;
        RECT 26.610 35.350 26.780 56.750 ;
        RECT 23.180 35.180 26.780 35.350 ;
        RECT 33.180 56.750 36.780 56.920 ;
        RECT 33.180 35.350 33.350 56.750 ;
        RECT 33.980 56.240 35.980 56.410 ;
        RECT 33.750 36.030 33.920 56.070 ;
        RECT 36.040 36.030 36.210 56.070 ;
        RECT 33.980 35.690 35.980 35.860 ;
        RECT 36.610 35.350 36.780 56.750 ;
        RECT 33.180 35.180 36.780 35.350 ;
        RECT 43.180 56.750 46.780 56.920 ;
        RECT 43.180 35.350 43.350 56.750 ;
        RECT 43.980 56.240 45.980 56.410 ;
        RECT 43.750 36.030 43.920 56.070 ;
        RECT 46.040 36.030 46.210 56.070 ;
        RECT 43.980 35.690 45.980 35.860 ;
        RECT 46.610 35.350 46.780 56.750 ;
        RECT 43.180 35.180 46.780 35.350 ;
        RECT 53.180 35.350 53.350 58.470 ;
        RECT 53.830 55.830 54.180 57.990 ;
        RECT 53.830 35.830 54.180 37.990 ;
        RECT 54.660 35.350 54.830 58.470 ;
        RECT 77.180 58.470 78.830 58.640 ;
        RECT 53.180 35.180 54.830 35.350 ;
        RECT 59.180 56.840 62.780 57.010 ;
        RECT 59.180 35.350 59.350 56.840 ;
        RECT 59.980 56.330 61.980 56.500 ;
        RECT 59.750 36.075 59.920 56.115 ;
        RECT 62.040 36.075 62.210 56.115 ;
        RECT 62.610 54.370 62.780 56.840 ;
        RECT 69.180 56.840 72.780 57.010 ;
        RECT 69.180 54.370 69.350 56.840 ;
        RECT 69.980 56.330 71.980 56.500 ;
        RECT 62.530 54.030 62.870 54.370 ;
        RECT 69.130 54.030 69.470 54.370 ;
        RECT 59.980 35.690 61.980 35.860 ;
        RECT 62.610 35.350 62.780 54.030 ;
        RECT 59.180 35.180 62.780 35.350 ;
        RECT 69.180 35.350 69.350 54.030 ;
        RECT 69.750 36.075 69.920 56.115 ;
        RECT 72.040 36.075 72.210 56.115 ;
        RECT 69.980 35.690 71.980 35.860 ;
        RECT 72.610 35.350 72.780 56.840 ;
        RECT 69.180 35.180 72.780 35.350 ;
        RECT 77.180 35.350 77.350 58.470 ;
        RECT 77.830 55.830 78.180 57.990 ;
        RECT 77.830 35.830 78.180 37.990 ;
        RECT 78.660 35.350 78.830 58.470 ;
        RECT 77.180 35.180 78.830 35.350 ;
        RECT 85.180 56.750 88.780 56.920 ;
        RECT 85.180 35.350 85.350 56.750 ;
        RECT 85.980 56.240 87.980 56.410 ;
        RECT 85.750 36.030 85.920 56.070 ;
        RECT 88.040 36.030 88.210 56.070 ;
        RECT 85.980 35.690 87.980 35.860 ;
        RECT 88.610 35.350 88.780 56.750 ;
        RECT 85.180 35.180 88.780 35.350 ;
        RECT 96.180 56.750 99.780 56.920 ;
        RECT 96.180 35.350 96.350 56.750 ;
        RECT 96.980 56.240 98.980 56.410 ;
        RECT 96.750 36.030 96.920 56.070 ;
        RECT 99.040 36.030 99.210 56.070 ;
        RECT 96.980 35.690 98.980 35.860 ;
        RECT 99.610 35.350 99.780 56.750 ;
        RECT 107.390 47.975 113.370 48.145 ;
        RECT 107.525 47.140 107.785 47.975 ;
        RECT 107.955 46.970 108.195 47.775 ;
        RECT 108.365 47.140 108.625 47.975 ;
        RECT 108.795 46.970 109.035 47.775 ;
        RECT 109.205 47.140 109.465 47.975 ;
        RECT 109.635 46.970 109.885 47.775 ;
        RECT 110.055 47.140 110.300 47.975 ;
        RECT 110.470 46.970 110.715 47.775 ;
        RECT 110.885 47.140 111.140 47.975 ;
        RECT 111.310 46.970 111.565 47.775 ;
        RECT 111.735 47.140 111.985 47.975 ;
        RECT 112.155 46.970 112.395 47.775 ;
        RECT 112.565 47.140 112.820 47.975 ;
        RECT 107.505 46.900 112.830 46.970 ;
        RECT 107.505 46.800 116.700 46.900 ;
        RECT 107.505 46.205 107.675 46.800 ;
        RECT 107.845 46.375 112.255 46.630 ;
        RECT 112.500 46.205 116.700 46.800 ;
        RECT 107.505 46.100 116.700 46.205 ;
        RECT 107.505 46.035 112.830 46.100 ;
        RECT 108.425 45.425 108.755 45.865 ;
        RECT 108.925 45.620 109.115 46.035 ;
        RECT 109.285 45.425 109.615 45.865 ;
        RECT 109.785 45.620 109.975 46.035 ;
        RECT 110.145 45.425 110.475 45.865 ;
        RECT 110.645 45.620 110.835 46.035 ;
        RECT 111.005 45.425 111.335 45.865 ;
        RECT 111.505 45.620 111.695 46.035 ;
        RECT 111.865 45.425 112.195 45.865 ;
        RECT 107.390 45.255 113.370 45.425 ;
        RECT 96.180 35.180 99.780 35.350 ;
      LAYER mcon ;
        RECT 19.910 57.915 20.100 59.900 ;
        RECT 19.910 35.920 20.100 37.905 ;
        RECT 24.060 56.240 25.900 56.410 ;
        RECT 23.750 36.110 23.920 55.990 ;
        RECT 26.040 36.110 26.210 55.990 ;
        RECT 24.060 35.690 25.900 35.860 ;
        RECT 34.060 56.240 35.900 56.410 ;
        RECT 33.750 36.110 33.920 55.990 ;
        RECT 36.040 36.110 36.210 55.990 ;
        RECT 34.060 35.690 35.900 35.860 ;
        RECT 44.060 56.240 45.900 56.410 ;
        RECT 43.750 36.110 43.920 55.990 ;
        RECT 46.040 36.110 46.210 55.990 ;
        RECT 44.060 35.690 45.900 35.860 ;
        RECT 53.910 55.915 54.100 57.900 ;
        RECT 53.910 35.920 54.100 37.905 ;
        RECT 60.060 56.330 61.900 56.500 ;
        RECT 59.750 36.155 59.920 56.035 ;
        RECT 62.040 36.155 62.210 56.035 ;
        RECT 70.060 56.330 71.900 56.500 ;
        RECT 62.530 54.030 62.870 54.370 ;
        RECT 69.130 54.030 69.470 54.370 ;
        RECT 60.060 35.690 61.900 35.860 ;
        RECT 69.750 36.155 69.920 56.035 ;
        RECT 72.040 36.155 72.210 56.035 ;
        RECT 70.060 35.690 71.900 35.860 ;
        RECT 77.910 55.915 78.100 57.900 ;
        RECT 77.910 35.920 78.100 37.905 ;
        RECT 86.060 56.240 87.900 56.410 ;
        RECT 85.750 36.110 85.920 55.990 ;
        RECT 88.040 36.110 88.210 55.990 ;
        RECT 86.060 35.690 87.900 35.860 ;
        RECT 97.060 56.240 98.900 56.410 ;
        RECT 96.750 36.110 96.920 55.990 ;
        RECT 99.040 36.110 99.210 55.990 ;
        RECT 97.060 35.690 98.900 35.860 ;
        RECT 107.535 47.975 107.705 48.145 ;
        RECT 107.995 47.975 108.165 48.145 ;
        RECT 108.455 47.975 108.625 48.145 ;
        RECT 108.915 47.975 109.085 48.145 ;
        RECT 109.375 47.975 109.545 48.145 ;
        RECT 109.835 47.975 110.005 48.145 ;
        RECT 110.295 47.975 110.465 48.145 ;
        RECT 110.755 47.975 110.925 48.145 ;
        RECT 111.215 47.975 111.385 48.145 ;
        RECT 111.675 47.975 111.845 48.145 ;
        RECT 112.135 47.975 112.305 48.145 ;
        RECT 112.595 47.975 112.765 48.145 ;
        RECT 113.055 47.975 113.225 48.145 ;
        RECT 110.815 46.415 110.985 46.585 ;
        RECT 115.930 46.130 116.670 46.870 ;
        RECT 107.535 45.255 107.705 45.425 ;
        RECT 107.995 45.255 108.165 45.425 ;
        RECT 108.455 45.255 108.625 45.425 ;
        RECT 108.915 45.255 109.085 45.425 ;
        RECT 109.375 45.255 109.545 45.425 ;
        RECT 109.835 45.255 110.005 45.425 ;
        RECT 110.295 45.255 110.465 45.425 ;
        RECT 110.755 45.255 110.925 45.425 ;
        RECT 111.215 45.255 111.385 45.425 ;
        RECT 111.675 45.255 111.845 45.425 ;
        RECT 112.135 45.255 112.305 45.425 ;
        RECT 112.595 45.255 112.765 45.425 ;
        RECT 113.055 45.255 113.225 45.425 ;
      LAYER met1 ;
        RECT 22.900 63.500 106.900 67.000 ;
        RECT 22.900 62.600 25.700 63.500 ;
        RECT 19.500 62.500 25.700 62.600 ;
        RECT 26.700 62.500 106.900 63.500 ;
        RECT 19.500 61.800 106.900 62.500 ;
        RECT 19.505 59.205 20.295 61.800 ;
        RECT 22.900 60.000 106.900 61.800 ;
        RECT 53.800 59.505 54.200 60.000 ;
        RECT 19.880 57.855 20.130 59.205 ;
        RECT 21.200 57.600 35.400 58.400 ;
        RECT 21.200 40.000 22.000 57.600 ;
        RECT 34.700 56.440 35.200 57.600 ;
        RECT 44.850 56.440 45.350 58.280 ;
        RECT 24.000 56.210 25.960 56.440 ;
        RECT 34.000 56.210 35.960 56.440 ;
        RECT 44.000 56.210 45.960 56.440 ;
        RECT 53.800 56.300 54.205 59.505 ;
        RECT 23.720 40.000 23.950 56.050 ;
        RECT 26.010 40.400 26.240 56.050 ;
        RECT 33.720 40.400 33.950 56.050 ;
        RECT 34.700 55.900 35.200 56.210 ;
        RECT 36.010 54.500 36.240 56.050 ;
        RECT 40.110 54.500 40.710 54.530 ;
        RECT 43.720 54.500 43.950 56.050 ;
        RECT 44.850 55.750 45.350 56.210 ;
        RECT 35.900 53.900 44.100 54.500 ;
        RECT 21.200 39.200 24.300 40.000 ;
        RECT 19.880 37.000 20.130 37.965 ;
        RECT 21.200 37.000 22.000 39.200 ;
        RECT 19.700 36.200 22.000 37.000 ;
        RECT 19.880 35.860 20.130 36.200 ;
        RECT 21.200 33.900 22.000 36.200 ;
        RECT 23.720 36.050 23.950 39.200 ;
        RECT 25.300 38.800 34.500 40.400 ;
        RECT 24.500 35.890 25.300 36.200 ;
        RECT 26.010 36.050 26.240 38.800 ;
        RECT 24.000 35.660 25.960 35.890 ;
        RECT 24.500 33.900 25.300 35.660 ;
        RECT 21.200 33.100 25.300 33.900 ;
        RECT 29.300 30.700 30.900 38.800 ;
        RECT 33.720 36.050 33.950 38.800 ;
        RECT 36.010 36.050 36.240 53.900 ;
        RECT 40.110 53.870 40.710 53.900 ;
        RECT 43.720 36.050 43.950 53.900 ;
        RECT 46.010 37.150 46.240 56.050 ;
        RECT 53.880 55.855 54.130 56.300 ;
        RECT 58.300 55.400 58.700 60.000 ;
        RECT 60.000 56.300 61.960 56.530 ;
        RECT 59.720 55.400 59.950 56.095 ;
        RECT 58.300 55.000 60.100 55.400 ;
        RECT 53.880 37.150 54.130 37.965 ;
        RECT 45.750 36.650 54.250 37.150 ;
        RECT 46.010 36.050 46.240 36.650 ;
        RECT 34.000 35.660 35.960 35.890 ;
        RECT 44.000 35.660 45.960 35.890 ;
        RECT 51.650 34.300 52.150 36.650 ;
        RECT 53.880 35.860 54.130 36.650 ;
        RECT 59.720 36.095 59.950 55.000 ;
        RECT 62.010 37.450 62.240 56.095 ;
        RECT 62.500 53.970 62.900 60.000 ;
        RECT 69.100 53.970 69.500 60.000 ;
        RECT 70.000 56.300 71.960 56.530 ;
        RECT 67.820 46.050 68.380 46.550 ;
        RECT 63.950 37.450 64.450 43.880 ;
        RECT 61.750 36.950 64.450 37.450 ;
        RECT 62.010 36.095 62.240 36.950 ;
        RECT 60.750 35.890 61.250 36.050 ;
        RECT 60.000 35.660 61.960 35.890 ;
        RECT 60.750 34.300 61.250 35.660 ;
        RECT 63.950 34.300 64.450 36.950 ;
        RECT 67.850 41.070 68.350 46.050 ;
        RECT 67.850 40.270 68.400 41.070 ;
        RECT 67.850 37.450 68.350 40.270 ;
        RECT 69.720 37.450 69.950 56.095 ;
        RECT 72.010 55.400 72.240 56.095 ;
        RECT 73.500 55.400 73.900 60.000 ;
        RECT 77.800 55.800 78.200 60.000 ;
        RECT 83.200 59.970 83.700 60.000 ;
        RECT 86.720 57.750 87.280 58.250 ;
        RECT 86.750 56.440 87.250 57.750 ;
        RECT 97.750 56.440 98.250 58.130 ;
        RECT 86.000 56.210 87.960 56.440 ;
        RECT 97.000 56.210 98.960 56.440 ;
        RECT 71.900 55.000 73.900 55.400 ;
        RECT 72.010 44.070 72.240 55.000 ;
        RECT 71.600 43.270 72.800 44.070 ;
        RECT 67.850 36.950 70.150 37.450 ;
        RECT 67.850 34.300 68.350 36.950 ;
        RECT 69.720 36.095 69.950 36.950 ;
        RECT 72.010 36.095 72.240 43.270 ;
        RECT 77.880 37.250 78.130 37.965 ;
        RECT 77.750 37.150 79.850 37.250 ;
        RECT 85.720 37.150 85.950 56.050 ;
        RECT 86.750 55.850 87.250 56.210 ;
        RECT 97.750 56.050 98.250 56.210 ;
        RECT 88.010 54.600 88.240 56.050 ;
        RECT 92.070 54.600 92.670 54.630 ;
        RECT 96.720 54.600 96.950 56.050 ;
        RECT 87.800 54.000 97.100 54.600 ;
        RECT 77.750 36.750 86.150 37.150 ;
        RECT 70.000 35.660 71.960 35.890 ;
        RECT 77.880 35.860 78.130 36.750 ;
        RECT 79.350 36.650 86.150 36.750 ;
        RECT 70.850 34.300 71.350 35.660 ;
        RECT 79.350 34.300 79.850 36.650 ;
        RECT 85.720 36.050 85.950 36.650 ;
        RECT 88.010 36.050 88.240 54.000 ;
        RECT 92.070 53.970 92.670 54.000 ;
        RECT 96.720 36.050 96.950 54.000 ;
        RECT 99.010 40.900 99.240 56.050 ;
        RECT 101.200 49.400 102.800 60.000 ;
        RECT 101.100 47.800 114.800 49.400 ;
        RECT 116.600 47.200 122.500 49.000 ;
        RECT 104.600 46.600 105.300 47.000 ;
        RECT 116.600 46.900 116.900 47.200 ;
        RECT 110.755 46.600 111.045 46.615 ;
        RECT 104.600 46.400 111.045 46.600 ;
        RECT 104.600 46.100 105.300 46.400 ;
        RECT 110.755 46.385 111.045 46.400 ;
        RECT 115.870 46.200 116.900 46.900 ;
        RECT 117.900 46.200 122.500 47.200 ;
        RECT 115.870 46.100 122.500 46.200 ;
        RECT 107.390 45.300 113.370 45.580 ;
        RECT 101.000 43.700 114.700 45.300 ;
        RECT 101.000 40.900 102.600 43.700 ;
        RECT 116.600 43.400 122.500 46.100 ;
        RECT 98.300 39.300 102.600 40.900 ;
        RECT 99.010 36.050 99.240 39.300 ;
        RECT 86.000 35.660 87.960 35.890 ;
        RECT 97.000 35.660 98.960 35.890 ;
        RECT 51.650 33.800 64.500 34.300 ;
        RECT 67.800 33.800 79.850 34.300 ;
        RECT 101.000 30.700 102.600 39.300 ;
        RECT 21.400 27.800 104.800 30.700 ;
        RECT 21.400 26.800 23.300 27.800 ;
        RECT 24.300 26.800 104.800 27.800 ;
        RECT 21.400 25.300 104.800 26.800 ;
      LAYER via ;
        RECT 34.700 57.600 35.200 58.100 ;
        RECT 44.850 57.750 45.350 58.250 ;
        RECT 40.110 53.900 40.710 54.500 ;
        RECT 67.850 46.050 68.350 46.550 ;
        RECT 63.950 43.350 64.450 43.850 ;
        RECT 86.750 57.750 87.250 58.250 ;
        RECT 97.750 57.600 98.250 58.100 ;
        RECT 92.070 54.000 92.670 54.600 ;
        RECT 104.650 46.250 105.150 46.750 ;
      LAYER met2 ;
        RECT 82.350 58.750 105.250 59.250 ;
        RECT 82.350 58.250 82.850 58.750 ;
        RECT 86.750 58.250 87.250 58.280 ;
        RECT 34.700 58.100 35.200 58.130 ;
        RECT 34.700 57.600 40.395 58.100 ;
        RECT 44.820 57.750 49.850 58.250 ;
        RECT 34.700 57.570 35.200 57.600 ;
        RECT 40.080 53.900 40.740 54.500 ;
        RECT 40.110 22.130 40.710 53.900 ;
        RECT 49.350 46.550 49.850 57.750 ;
        RECT 82.350 57.750 87.250 58.250 ;
        RECT 91.475 58.100 91.925 58.120 ;
        RECT 67.850 46.550 68.350 46.580 ;
        RECT 49.350 46.050 68.350 46.550 ;
        RECT 67.850 46.020 68.350 46.050 ;
        RECT 82.350 43.850 82.850 57.750 ;
        RECT 86.750 57.720 87.250 57.750 ;
        RECT 91.450 57.600 98.390 58.100 ;
        RECT 91.475 57.580 91.925 57.600 ;
        RECT 104.750 57.090 105.250 58.750 ;
        RECT 104.650 55.750 105.250 57.090 ;
        RECT 92.040 54.000 92.700 54.600 ;
        RECT 63.920 43.350 82.850 43.850 ;
        RECT 40.110 21.530 44.305 22.130 ;
        RECT 92.070 21.150 92.670 54.000 ;
        RECT 104.650 46.220 105.150 55.750 ;
        RECT 92.025 20.550 92.715 21.150 ;
      LAYER via2 ;
        RECT 39.850 57.600 40.350 58.100 ;
        RECT 91.475 57.625 91.925 58.075 ;
        RECT 43.660 21.530 44.260 22.130 ;
        RECT 92.070 20.550 92.670 21.150 ;
      LAYER met3 ;
        RECT 39.825 58.100 40.375 58.125 ;
        RECT 39.825 57.600 91.950 58.100 ;
        RECT 39.825 57.575 40.375 57.600 ;
        RECT 43.635 22.130 44.285 22.155 ;
        RECT 43.635 21.530 45.860 22.130 ;
        RECT 43.635 21.505 44.285 21.530 ;
        RECT 92.045 21.150 92.695 21.175 ;
        RECT 88.010 20.550 92.695 21.150 ;
        RECT 92.045 20.525 92.695 20.550 ;
        RECT 33.400 -11.060 65.260 19.340 ;
        RECT 69.780 -10.480 101.640 19.920 ;
        RECT 33.400 -42.660 65.260 -12.260 ;
        RECT 69.780 -42.080 101.640 -11.680 ;
        RECT 33.400 -74.260 65.260 -43.860 ;
        RECT 69.780 -73.680 101.640 -43.280 ;
        RECT 33.400 -105.860 65.260 -75.460 ;
        RECT 69.780 -105.280 101.640 -74.880 ;
        RECT 33.400 -137.460 65.260 -107.060 ;
        RECT 69.780 -136.880 101.640 -106.480 ;
      LAYER via3 ;
        RECT 45.230 21.530 45.830 22.130 ;
        RECT 88.040 20.550 88.640 21.150 ;
        RECT 64.840 -10.920 65.160 19.200 ;
        RECT 101.220 -10.340 101.540 19.780 ;
        RECT 64.840 -42.520 65.160 -12.400 ;
        RECT 101.220 -41.940 101.540 -11.820 ;
        RECT 64.840 -74.120 65.160 -44.000 ;
        RECT 101.220 -73.540 101.540 -43.420 ;
        RECT 64.840 -105.720 65.160 -75.600 ;
        RECT 101.220 -105.140 101.540 -75.020 ;
        RECT 64.840 -137.320 65.160 -107.200 ;
        RECT 101.220 -136.740 101.540 -106.620 ;
      LAYER met4 ;
        RECT 45.225 22.130 45.835 22.135 ;
        RECT 48.340 22.130 101.650 22.200 ;
        RECT 45.225 21.680 101.650 22.130 ;
        RECT 45.225 21.530 49.170 21.680 ;
        RECT 45.225 21.525 45.835 21.530 ;
        RECT 48.340 18.945 48.860 21.530 ;
        RECT 88.035 21.150 88.645 21.155 ;
        RECT 83.290 21.130 88.645 21.150 ;
        RECT 64.660 20.610 88.645 21.130 ;
        RECT 64.660 19.940 65.180 20.610 ;
        RECT 83.290 20.550 88.645 20.610 ;
        RECT 33.795 -10.665 63.405 18.945 ;
        RECT 64.660 14.670 65.260 19.940 ;
        RECT 84.720 19.525 85.240 20.550 ;
        RECT 88.035 20.545 88.645 20.550 ;
        RECT 101.130 20.520 101.650 21.680 ;
        RECT 48.340 -12.655 48.860 -10.665 ;
        RECT 33.795 -42.265 63.405 -12.655 ;
        RECT 48.340 -44.255 48.860 -42.265 ;
        RECT 33.795 -73.865 63.405 -44.255 ;
        RECT 48.340 -75.855 48.860 -73.865 ;
        RECT 33.795 -105.465 63.405 -75.855 ;
        RECT 48.340 -107.455 48.860 -105.465 ;
        RECT 33.795 -137.065 63.405 -107.455 ;
        RECT 48.340 -138.060 48.860 -137.065 ;
        RECT 64.740 -138.060 65.260 14.670 ;
        RECT 70.175 -10.085 99.785 19.525 ;
        RECT 101.120 14.060 101.650 20.520 ;
        RECT 84.720 -12.075 85.240 -10.085 ;
        RECT 70.175 -41.685 99.785 -12.075 ;
        RECT 84.720 -43.675 85.240 -41.685 ;
        RECT 70.175 -73.285 99.785 -43.675 ;
        RECT 84.720 -75.275 85.240 -73.285 ;
        RECT 70.175 -104.885 99.785 -75.275 ;
        RECT 84.720 -106.875 85.240 -104.885 ;
        RECT 70.175 -136.485 99.785 -106.875 ;
        RECT 84.720 -137.480 85.240 -136.485 ;
        RECT 101.120 -137.480 101.640 14.060 ;
  END
END osc
END LIBRARY

