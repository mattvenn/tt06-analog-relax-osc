magic
tech sky130A
magscale 1 2
timestamp 1710835479
<< psubdiff >>
rect 21282 6460 21306 7326
rect 22216 6460 22240 7326
<< psubdiffcont >>
rect 21306 6460 22216 7326
<< locali >>
rect 22500 9374 23340 9380
rect 21800 9317 22200 9320
rect 21800 9283 22163 9317
rect 22197 9283 22200 9317
rect 21800 9280 22200 9283
rect 22500 9226 23186 9374
rect 23334 9226 23340 9374
rect 22500 9220 23340 9226
rect 21290 6460 21306 7326
rect 22216 6460 22232 7326
<< viali >>
rect 12506 10806 12574 10874
rect 13826 10806 13894 10874
rect 22163 9283 22197 9317
rect 23186 9226 23334 9374
<< metal1 >>
rect 4580 12520 21380 13400
rect 3900 12360 21380 12520
rect 3901 11841 4059 12360
rect 4580 12000 21380 12360
rect 10760 11901 10840 12000
rect 4240 11620 7080 11680
rect 4240 11520 6940 11620
rect 7040 11520 7080 11620
rect 8970 11650 9070 11656
rect 4240 8000 4400 11520
rect 6940 11180 7040 11520
rect 8970 11150 9070 11550
rect 10760 11260 10841 11901
rect 11660 11080 11740 12000
rect 11660 11000 12020 11080
rect 8022 10900 8142 10906
rect 7180 10780 8022 10900
rect 8142 10780 8820 10900
rect 12500 10874 12580 12000
rect 12500 10806 12506 10874
rect 12574 10806 12580 10874
rect 12500 10794 12580 10806
rect 13820 10874 13900 12000
rect 14700 11080 14780 12000
rect 15560 11160 15640 12000
rect 16640 11994 16740 12000
rect 17344 11550 17350 11650
rect 17450 11550 17456 11650
rect 19550 11620 19650 11626
rect 17350 11170 17450 11550
rect 19550 11210 19650 11520
rect 14380 11000 14780 11080
rect 18414 10920 18534 10926
rect 13820 10806 13826 10874
rect 13894 10806 13900 10874
rect 13820 10794 13900 10806
rect 17560 10800 18414 10920
rect 18534 10800 19420 10920
rect 18414 10794 18534 10800
rect 8022 10774 8142 10780
rect 20240 9880 20560 12000
rect 20220 9560 22960 9880
rect 20920 9350 21060 9400
rect 23320 9380 24500 9800
rect 13564 9210 13570 9310
rect 13670 9210 13676 9310
rect 20920 9250 20930 9350
rect 21030 9320 21060 9350
rect 23174 9374 24500 9380
rect 22151 9320 22209 9323
rect 21030 9317 22209 9320
rect 21030 9283 22163 9317
rect 22197 9283 22209 9317
rect 21030 9280 22209 9283
rect 21030 9250 21060 9280
rect 22151 9277 22209 9280
rect 20920 9220 21060 9250
rect 23174 9226 23186 9374
rect 23334 9226 24500 9374
rect 23174 9220 24500 9226
rect 12790 8770 12890 8776
rect 4240 7840 4860 8000
rect 4240 7400 4400 7840
rect 5060 7760 6900 8080
rect 3940 7240 4400 7400
rect 4240 6780 4400 7240
rect 4900 6780 5060 7240
rect 4240 6620 5060 6780
rect 5860 6140 6180 7760
rect 12790 7490 12890 8670
rect 9150 7330 10850 7430
rect 12350 7390 12890 7490
rect 10330 6860 10430 7330
rect 12150 6860 12250 7210
rect 12790 6860 12890 7390
rect 13570 8214 13670 9210
rect 14320 8654 14560 8814
rect 20200 8740 22940 9060
rect 13570 8054 13680 8214
rect 20200 8180 20520 8740
rect 23320 8680 24500 9220
rect 13570 7490 13670 8054
rect 19660 7860 20520 8180
rect 13570 7390 14030 7490
rect 15550 7430 15970 7450
rect 13570 6860 13670 7390
rect 15550 7350 17230 7430
rect 15870 7330 17230 7350
rect 14170 6860 14270 7160
rect 15870 6860 15970 7330
rect 10330 6760 12900 6860
rect 13560 6760 15970 6860
rect 20200 6140 20520 7860
rect 21254 6140 22334 7462
rect 4280 5060 22334 6140
<< via1 >>
rect 6940 11520 7040 11620
rect 8970 11550 9070 11650
rect 8022 10780 8142 10900
rect 17350 11550 17450 11650
rect 19550 11520 19650 11620
rect 18414 10800 18534 10920
rect 13570 9210 13670 9310
rect 20930 9250 21030 9350
rect 12790 8670 12890 8770
<< metal2 >>
rect 16470 11750 21050 11850
rect 16470 11650 16570 11750
rect 17350 11650 17450 11656
rect 6940 11620 7040 11626
rect 7040 11520 7970 11620
rect 8070 11520 8079 11620
rect 8964 11550 8970 11650
rect 9070 11550 9970 11650
rect 6940 11514 7040 11520
rect 8016 10780 8022 10900
rect 8142 10780 8148 10900
rect 8022 4426 8142 10780
rect 9870 9310 9970 11550
rect 16470 11550 17350 11650
rect 18295 11620 18385 11624
rect 13570 9310 13670 9316
rect 9870 9210 13570 9310
rect 13570 9204 13670 9210
rect 16470 8770 16570 11550
rect 17350 11544 17450 11550
rect 18290 11615 19550 11620
rect 18290 11525 18295 11615
rect 18385 11525 19550 11615
rect 18290 11520 19550 11525
rect 19650 11520 19678 11620
rect 18295 11516 18385 11520
rect 20950 11418 21050 11750
rect 20930 11150 21050 11418
rect 18408 10800 18414 10920
rect 18534 10800 18540 10920
rect 12784 8670 12790 8770
rect 12890 8670 16570 8770
rect 8022 4306 8732 4426
rect 8852 4306 8861 4426
rect 18414 4230 18534 10800
rect 20930 9350 21030 11150
rect 20930 9244 21030 9250
rect 18405 4110 18414 4230
rect 18534 4110 18543 4230
<< via2 >>
rect 7970 11520 8070 11620
rect 18295 11525 18385 11615
rect 8732 4306 8852 4426
rect 18414 4110 18534 4230
<< metal3 >>
rect 7965 11620 8075 11625
rect 7965 11520 7970 11620
rect 8070 11615 18390 11620
rect 8070 11525 18295 11615
rect 18385 11525 18390 11615
rect 8070 11520 18390 11525
rect 7965 11515 8075 11520
rect 8727 4426 8857 4431
rect 8727 4306 8732 4426
rect 8852 4306 9046 4426
rect 9166 4306 9172 4426
rect 8727 4301 8857 4306
rect 18409 4230 18539 4235
rect 17602 4110 17608 4230
rect 17728 4110 18414 4230
rect 18534 4110 18539 4230
rect 18409 4105 18539 4110
<< via3 >>
rect 9046 4306 9166 4426
rect 17608 4110 17728 4230
<< metal4 >>
rect 9045 4426 9167 4427
rect 9668 4426 20330 4440
rect 9045 4306 9046 4426
rect 9166 4336 20330 4426
rect 9166 4306 9834 4336
rect 9045 4305 9167 4306
rect 9668 3884 9772 4306
rect 17607 4230 17729 4231
rect 16658 4226 17608 4230
rect 12932 4122 17608 4226
rect 12932 2934 13036 4122
rect 16658 4110 17608 4122
rect 17728 4110 17729 4230
rect 16944 4000 17048 4110
rect 17607 4109 17729 4110
rect 20226 2812 20330 4336
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0
timestamp 1685868990
transform 1 0 21314 0 1 9070
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_8  x1 ~/.volare/volare/sky130/versions/78b7bc32ddb4b6f14f76883c2e2dc5b5de9d1cbc/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 21478 0 1 9068
box -38 -48 1234 592
use sky130_fd_pr__cap_mim_m3_1_39BNLG  XC1
timestamp 1710760421
transform 1 0 9866 0 1 -11812
box -3186 -15800 3186 15800
use sky130_fd_pr__cap_mim_m3_1_39BNLG  XC2
timestamp 1710760421
transform 1 0 17142 0 1 -11696
box -3186 -15800 3186 15800
use sky130_fd_pr__nfet_01v8_L9BG78  XM1
timestamp 1710760421
transform 1 0 8996 0 1 9210
box -396 -2210 396 2210
use sky130_fd_pr__nfet_01v8_L9BG78  XM2
timestamp 1710760421
transform 1 0 17396 0 1 9210
box -396 -2210 396 2210
use sky130_fd_pr__pfet_01v8_5Q5MA6  XM3
timestamp 1710760421
transform 1 0 14196 0 1 9219
box -396 -2219 396 2219
use sky130_fd_pr__pfet_01v8_5Q5MA6  XM4
timestamp 1710760421
transform 1 0 12196 0 1 9219
box -396 -2219 396 2219
use sky130_fd_pr__nfet_01v8_L9BG78  XM5
timestamp 1710760421
transform 1 0 4996 0 1 9210
box -396 -2210 396 2210
use sky130_fd_pr__nfet_01v8_L9BG78  XM6
timestamp 1710760421
transform 1 0 6996 0 1 9210
box -396 -2210 396 2210
use sky130_fd_pr__nfet_01v8_L9BG78  XM8
timestamp 1710760421
transform 1 0 19596 0 1 9210
box -396 -2210 396 2210
use sky130_fd_pr__res_high_po_0p35_NFQ4JE  XR1
timestamp 1710760421
transform 1 0 10801 0 1 9382
box -201 -2382 201 2382
use sky130_fd_pr__res_high_po_0p35_NFQ4JE  XR2
timestamp 1710760421
transform 1 0 15601 0 1 9382
box -201 -2382 201 2382
use sky130_fd_pr__res_high_po_0p35_QPS5FG  XR3
timestamp 1710760421
transform 1 0 4001 0 1 9582
box -201 -2582 201 2582
<< labels >>
flabel metal1 5140 12500 5340 12700 0 FreeSans 256 0 0 0 VDD
port 1 nsew
flabel metal1 4660 5360 4860 5560 0 FreeSans 256 0 0 0 VSS
port 2 nsew
flabel metal1 23380 9240 23580 9440 0 FreeSans 256 0 0 0 osc_out
port 0 nsew
flabel metal1 12790 6760 12890 8670 0 FreeSans 1600 0 0 0 osc_a
flabel metal1 13570 6760 13670 9210 0 FreeSans 1600 0 0 0 osc_b
flabel metal2 8022 4306 8142 10780 0 FreeSans 1600 0 0 0 left_cap
flabel metal2 18414 4230 18534 10800 0 FreeSans 1600 0 0 0 right_cap
flabel metal1 4240 11520 6940 11680 0 FreeSans 1600 0 0 0 cset
<< end >>
